--
--Written by GowinSynthesis
--Product Version "V1.9.8.11 Education"
--Mon Jul 24 09:51:06 2023

--Source file index table:
--file0 "\/home/cod3r/Data/Gowin/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\/home/cod3r/Data/Gowin/IDE/ipcore/DVI_TX/data/rgb2dvi.vp"
`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
n9djzkmMiau/ZFbYlXd99E90bX+ysAJqTLVkQsG6tiUrKJJ0KuA5B81N+Fk+S7oTwc7H3Z9CLi3D
zJhqJB+Cy3jN1Efn8oS2VvxaYEwBU4yAuanYK5EEsaPSOpLprxecR5TPSBAyvbt8vAgmfdXB2Cce
MZYajlZR8WEYMPSKwOsfQZ1dkS0UyQorMfyeVpwpu7959FXG1+IR8FtOOCgFxYgXyL8aaQKaor0h
Mmgr2/3+TUvS/0kHjKUmaXo8EUCSsOOqj88pKwQV37pf5xHhS/H7pUbD5e7nUxOQpsyDhIX5GOpW
/xUmSAf46198FG3fKlZh5ncJobjC8brf17gAWQ==

`protect encoding=(enctype="base64", line_length=76, bytes=69408)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
4ZMXj6xgWHkyWJmXTPGaiQaw3POCHn4vhXncg91PzPx7MClbiPMsTLSJGAz1HwFqI5F4F4a8zmor
raBVxaiAtrbGIduPRHSaneSahk3tXUT3/gvH59S9KfAfRR77b5vCh0uv8S9+V8FKL94EDVyg1cV6
zB74rVzq98w5E3bhnx3TdZbL/29SOrB7gc3gOQvwOZChpUjw1CwiFa5n3J5+oCQHjT7+I1ACSZBM
vYUFr7evvKssgs+8fQERRWNcTOuezNWND0rz+6DLnMMwbXXS3owSbkkOVZm0HmmrbSm3FZHpipM8
1DSZ+0QExvkK4zw4fet4ujCrhLoakQdQS8cd6m8+cPFqrzPPRwYvdmJd9E+DjXqF9SvRQPvCpj6v
++gYetaXUtH4diovPbBU8Uy2Hzy4U0GBsw2PjeEwUtMBwZ0eMgrD1Id8ISOOJUPGwK/HtKjh7H4n
PCuOHLERS3M8lPSSGj1rJ9Eg1pfzOOVUv545EdCqS0UQX+6UXTCGedjRDIfNA/AF3SXLQJybQK/V
dEcyKRUqZUg0X73efCN5eZK9PMbo0J3gmPs9xID4SitUGfcEmVBRdAMH4Oc1SzF9ITDhcL444s/8
IGa84eWRMFwd8RJoz7Tnf/sRpTfcxS9dhWqw+COAd3IH7jh9vRZVVQlvWG1XnyuG74W6V/9doxp5
bQAyHU3We3EBT6KXtB0AFesXbjQ9sEbqbNbjHCFab3Wegv1YUoE3SbaXMPvwDkksXvVn/dBYsu6l
rI4c1psXFMp2UYYXfxPZmA4oaXljn8JlxAyUOL7XFeYxAB+L3kFX/HYvHNBsePf7in2TvJvWaWv/
4hUa8znjwq6dcucfulZa1wOpxukI1gp4xRpXtlZk6xagQw7r6qc6FxY2WKoijPK74UFmQPyRXQRa
1FEPcJNTCmMAV6dH0vi5g5C7N/IJ85VuPdF8URfjf1aQU/4/3CEZq6zCfMvEsrUAWHS8b38CYDef
jQ0vsNttlBEhY7/dXxPZHmb+ByezNe/lWF2Q0ubq8iYhNEQYpz2JMk+sgTTzzIrYntN0AVzdCyXU
wCLTRFXG223CiYCGDysugb2WoI/umIAdEaA65gT7FE9N6VSOcPmhPH2pinCmpXLIWMB//m79GzZG
9ptF3vnNMGJVF72W2nH9MxP05hYFHNaTcqkkHKY7IBUsSLPEq7ad7zO/bgU2diDRyZeSG1ks4sWu
cgrEN7ReqXy2JLMNosb0HFo/SB0IJyUfDjJhDXUmv4lYomJQX9qehx36QgvQmSD6veQU0HlcFNCS
kZ2Vk//US1raYt3WiT8DVFxCmsOJFfGEqQ0FWvX/w8paGioFWHac3ohHYr/YnFeIfA8aM0JaOMRf
XjIH0BzHUd6clcpVzrRSpvAP1qW8s5IcmipQl/jV3iYMisn05u5JrMcIGEPhG1p1abFpm83MlFtt
+jeYkd7I+7v23uz+e9PUOBbSbezxq57MsSxuMU3kCtKLaint2IOwnhGmgPMaVxefgEDSMVP92wqU
HW9RIoiRb/uNM7k1UTL0gwdhDPGIzanax0ZFDlDWHA7VJaKb3IKe+H6GY/gi4skDB39cO97OlCyb
pJIb1ns8z71iEX2gHaOChtud9pw/VyzOB9EtOnFSKar7isqmBpNFS0N43zpJeBUTt2hmc1EJI4kW
Srqa/FYMrJ76+VBp/YYRkNHBLZiFDpWtoWi2asqWHE/NWrk3z/PnLpKWv55ER1mZ6H1zQ63Qsj8q
oBeh8Ivrh/fWqlpqgED4P7u3vkFEDJ4t8rx6kzCDCaAF7LzhNBs+C0b3WaPn0oPxb8yQLA+eQ+/q
sjiNQ86gIPu6Bh7HLQgXZz2ADqlDZ0gtHCCl2kjDYEyReSYHWrHBF+0M5KkXIQzuKp4U0G5mtH2z
x1TNy21M9SzRAleszOIE8bS3G3Qgu9n7LoTsI83lgABqFmYxwhymg47mZY65NuWpeUwykPP2MfHC
bTPnHOZOhpvsSCquIYpDST6Fo8V7NopQ+JM/s17+1+10wPnznDqGi+8S7sn27beeCp6zm/8nn215
yXLF8N+PY/jPCIhnDKNyezRpFDEmVIME/DhDLs+sFeXhI4KKwrGP/qEmT3NshOPS93gnhqliTOFi
oaVFR88cvwGfFWqL7Y59XJykHqODO8lA8x0b4fwUMu4AAE4IJ879FTPvbpranIB27JyinTB1Ic/y
bLDv0+1L6erCFV9j9yfIpfOQHeWE+Etgh7bMdkBw5mi+Bx+CA2WrQouAIfH79p/d0X0vVaCaZ1FF
oOeAGANoZ4u6A3Q7pzwiNyALU9g1ta8lhhPMf6NFPhsMOUfn8GzNSO1GSpznWHvMcldyhSA/4shL
IOylVb9RjbYicVZJMyJIGN5AO81HzWgtjxfar8LjsEjAvBxVAgEypJkHo1HsBjMg0ZZiPYgO1yHZ
X03sHMBPwAKi+dTMlXmLAX1h5tnq8HHi3ZPk4xzoAdVrSKpMo1oBNO3/ToizODx4PlT3Ka5sja8+
wrRuZEnO+s1gtVF3u1eZk9esffKOTz7QklI+2AipybdQlh9/mbMd9RPnmrNadY1NUTOoMYLF6kut
vBV8qPHvMNxBs+6zXfoo2WGyQnKR5dJoiIs3fAV0CH2OhzjhJ/IvO0QD5MhthaW5UVyovk3XTDES
aZsLmV/5VFYdV7+4YAvoQS+1wKbHaR9PkCsonZUwUnS+g2547ARXysERJSJT0HKC6/nggUa7nUG9
kz21qXVlzxL8I7ojt6VGDXgFkSgoD9/Gp+LssOdr4A2xkTKvY3GHfPoZr/tp1OPtHLSPgyDCIjfN
cKWflkMJnLAJKZ67IEGSl1bkB1yWKnHK4JEYYuVLJiP/O+7aibVl8jf+eQTef2XLUOsxWj9NYQWE
qGsEtIyymPIvtkUnY51Z0Oh9njSMcmHN0LSCk5yTiYzXTD/SpWDdBjNF66BTVb6xM4dIK0OSNsCD
mu1gHsrvUm0Q7YuB6E7wmXxCv6EmobK/1mxN6RTB3P1MyvmZUBu6ZOp6uEnMSPRLKMkbsGML+jvo
AkJiZyfZkLFo+dG1E0l59IvYVBMiSveQTBccLDmN+lol3v3uLFhUG3ylqQbQ7/en0x0xSrPMYQEK
+vLepsFNW/GHSvkBGIJ1UCj8QcOLgMilAHCY2rLZ4o7nP30GL6ievhObGdJmtnEs29xKd0LGvDKh
AGkL7pc0Z3on2suwBV8O+j1pvvJCw3DYqUSWyB46bzd+fFpk3YUKxwwcYalz4VzExxoRBXsbeqI9
FbqQw1fxMkZjaJ/924sB6r1XsQYgyTN6dRXqCZUrufgSYV14+FflPnEiVxIGWLRRO2Cd0fYFeNCM
JwIYfKpGWXKzKN1B2pmBXyXHYzSluJ/lGMlUdU6YYjcTrOK1AQLqQhQ+SX3xONyWTAeon1PTu7w9
wnF8lNNwqOV4o7th25FI/Ws9Cxw6x/XfqXJVqAp9wU4cUex+zCeEClbafxAzXJrZAleenxB4Uvou
35qVTExdgv6NcEXIo4l8GWSgxnsB2v+apJSrJCQoUkwtfXNU8AqdIlkdyqI8WNyhmE1xrZ3NyRwU
OePayxLgS6Yen7e/bNEkXaeISOydQq1HbzHeuvnLQqmTHp/Eq9kGJJxBFdsTdpx5YOjZjHlyPCmS
Zp78wSeciQwq48JsBpuFma/9e8qng3tNFjqKZLwpaI1h1bp27jwQA0EjFxD6QprEdK6a3G4BuHLW
609kWNPPJyNsER/4TfP0ZS2wid9H1ZreAzQNn0l4An1gszn1lE+CYQECQyMiHDyQY9iERjF243IU
ttN56kxcaMJaL+88v36I1+nOqaskMdVurz6z0x/TLPqZ4FBnErDVb6YCqTugXZyn1fPCQ/1U/v8I
e/Q3tjq5f3nESr72HVdPOpFlS/ADL2Wgz7aXcuPXSAYyNeMpzZ3mvpVNXMkKA3kRxtOhN5LFoBP6
KPtNGZ+dlcE5aOoq67m/ndRyKEbeZO7GLbWWd52YrLiYm6oA6DDgDdvj3JrtFkQKyGSt0wgnG69x
uaFykRmot6lmi3UBBCoJovSXlYyPI1zUN8dizhxJRImF9N73MGhDYCGoMBfZ+oqcxzT/FVwESE1u
cfj1bMCCv9mBmMGtFck8MiK8Gnw08nimEQaksBz60EYz3cbIbMNwOiJu8vuo6f6LFIPpgZCVODLq
d1wOFU52GCajO58L9DWTuz+1puGMClW4cA9Zhi/i1uqyh5fS71YpEHO2f6LZOjbVl5pooj3rXumt
JlT//4oo4bEkS0XxAzZGpArRFXeYs0Y8/IrzJv3o0RUiZsoenElu3ORMrKhzGSGKN99k+FZ02Kwi
19Q/UPAAnjERBXhsGKCmQTXuov1oRAElr8y3IrRiaoQCVFuqnEtTgp/o+SuOQU7sCWDeLPq3vWto
PTXPUHiX5sMPehErYUrf3HI4XW7X2jGAcYuBNJUOf/GvXdmCpmqZDDGQ2M1g3/sZeNJpnv1ZPUrg
ss52FTOcTQ+CvHnwyiWluNYadoZudR5s0VKSupmIM205IDC8FusHW0D1vS5TFFXCVg/hml0mACEi
yhnXmpcpGwGzsZuuLZqmmYOL8gmSDvCNYc+QaDqspqGVioDkmgbkI4qNUugsnpInbCEfX8GagTVE
1G/9Ee4zvjsePLsFCsie0ZxsEitCrngKyI3MHGVVDA4311/0/eJpVtJR5B8KPPPcwMpdoD3DPOY0
llbU38uTGgswFft+BV4/2wXYi9sNLZYUpCyorohYyfx96S9iU+InR8u22g/HKHKqtCcJ6pqRtLXc
6D2s1gGyZ9vEscnvHrGn9N28UBMo/KVTxQ7mS90f3BKWyqcBK7OtLPaMk6Wf1/KeNSLbqx5lIadF
iTbH7iZKu5KpwSjusgL1ugVlWkHaiQn7SFlvvhlO1Rlp1+87NAyrj1KsshwvbgJT58QRA9zcZbch
yT4uvIBzTiGUYSwLmK3FcWzImM3e+q54tRj5+zWoOUD7ZcofbZZDa0Cwzuf1szwP85DR1Vcwbmle
+VDekGKZjYQvgJH/Yn950ly+31f2FVthiqqbhROsGl9NOpr0xRVe1TRLJr467wO2f70bRAnXSmLO
ZIUG9HmWabNUy8vTqpmXtuscVK0Go4F3E7jUy6bzlwvpNNEsX6iL7/nqGzb+0Am2mi0kS5MbhHAb
e6aRD6BgXzhPbPUITbm+DJMSRfSjF0jGHBgVZ0CU8BRB64iTzkztfYEU4aVl8PPKmtcse4IkDhMo
seooONtEO6xkaBrUqa1JlaOPx91+BaT7sNA3xYg9iOwI1egA+ZSQrakjGa5dk/KGyb0Bs+zVfNAe
SzE+31MPA3FYyzZdB5wVFDihnRKJjVzKSP5pbPjLInYV2FVwTuRB3dC10idwmnKdq6wUhfb6AFJ9
fZEcNQ69YQzCG9+9YSkoFTTXvdWFlEzbi9gr4GmodwpdsoKRg4XoxcAoTDLizEI21rRnuCFAZEcD
2yHSrCqX+HbcCmwxfvjfUDGjjxLwAJ9Wqwmc8dEvTwuPB+Lm4cXnvEN4PtvS6uvEQxOSkVMKDLUw
TED0DQo/ZwQe59hA6R3qDHB0om5WnQltFfB04fzPA7/GvLOLZ9JFbNwK3000V4Od3/JKnKVykbLl
LMeXoG6DJO7NKUKhiu0MG44d+ZEN1sfFkwrkTe3/yY/ppDgtVanw+louV/k9DWvjGFY0bdg5iAhr
/9fPXkg878F7iGFC+Pxi/EQ6fyVMOg7HumOyKRSYNBUMT0SE+olQGV5BNsNlK7smSZwVY9HXm8nI
KuIsTZclJsDAG8HMkPzFzvqe37uDLHJIh9zQWR44XjzY11tJDNsLaFVJwZ3iWsRGEKwh2exRV2m5
H2f3E1VaWEsuGyPjUx7z6puNzEfI7fEUZOauaSGSJXkDlASK+Cqb0PjO5Jx6g0LlrkWYm7z5ygJw
3ImyVXXKxCBqvKnpvEsJcxiPiyuBUlmzCkCOLhF1bAMZR7j/Lq7R0TVFZ1pRhV8LewR70xMgDVPk
3SLQePM6DutBPcOT7aG6f9Ni7tAN1PEv2sdhf7owotCvr32Seyghgrzys/7NgZXzTkzR0Wx2O3ZV
8vdhMjjsCLT2MZTNBzyWcPMNhSzKkAFXGdQVbH8G7ZAEFh1fihS1pTE09g5ZdBxWA8WuWxtRVOIC
a+JXNoQWWDl+r5+Vt4mjzV06Nf0tONRrtTLAbtKhRzzK7Hflyuw14Lj+NeKbhhlJ5/ifvgyfigH9
AmfcOA4vb2NI/2eGhwFePdv3c26BEjx5EMZYCJTqkS+zEWrWphzzp/gft4mEys6MspE0F2xOVyAA
cnxZF2iiYhnFXDg0jzl5EQjuUFbqh4NxToMasTXKFW5f4+vqtcIm5INLVb8ahyjgl9k/vnXdY+HT
ssqHPUpcImeeNSd5om5SFRYEnehqL4b0ep+TW8VRTySyeVonawdeoxrj04u1cocKbl7bBmcD4Aei
4lCdCzZytiHEky9SY6ZNCn/br1hQCpnRNunVPGHO5AujYEvMP+4jEnlA90+ncaCT6opoDGoLKUMk
YN+bya7F1wm/tm00nyI78rhjFCqFnEoEDWB5SqvEOqZf0FX+EbfmdO9LgWCSfNpYj1RwvrY7hHyd
ZxpeqyPEiAwUcCLPxVfB/N6AdB7mJLUCuemXajS3ASMCX0RpOBiFgGzFPupdb3KY/R1vMhHufxs/
WGMM+TXB2gklj+OQrDOEAoO2ya/eVanWL1Q4Cx/nXDdNS9PsFYngep7l6dqwY10L5qe/sst/KVHL
QgmyXkHwqftEwebUqLRMZP8LSJpPWlFliUTl6OJsIATczgO4m4RScJGgUwUVcUjgMnfKpTmnp6/c
NuqCH46LSlRYsCYUktCwYfHtcSPq3VkRDJ4OckqRvUPbhfq3n1sfMPv+w20sIAR8V4EmR45E7V0B
TZoHHJM7R9jwilAMS5XVQHeQBINFTf/glzeH04N52OimYPK1N6VACaQj/BLuzxs4m6sHy5/L6U3r
FVLk0ETRknjkWOFYU6mrlNR21Koogj99QhGB9UTrwDIMWqy3ehr3gRKoh546xJNuT/dWhUh15AXK
eqNianFR4yhwk9R1zPSyr/vdpkiQpcKJqtZhjrZdkH8HIDH45IZJEkRubjEXpz6QWcPoCYWt/TWi
jy5Z2xDZaXrDyBqiLL/9p/HbsjkITmJ0LqfyfWPQB3/z8j9f+Fzx30sJXg5gRcXjamcNeT9d5UJm
3Av0eDs7qpZxpP7VHN1Kw212mZ4VJC/lCllz+FriDlVNlwGdYep/5ObgRROyokXxmOA7zFW+JBNJ
ceuxayHBen6rGcQTuU7g1wcIZ4JCV4Xb43YDNh2/jN0tz4bDeFhcHyc572+6zINEL8flejEI1qdf
sGIoOfWsQEAUJcTRLcF1/ph8yVGrFtb+2cD5UqPB7gBg9WtQcla5aBhucaa4qytySY477kAYBedB
zkSh+eej8g5iE4a65e9LW17rX4ajLEv/w5a40aSGBDZTuU3tGCTj2BybdyTnUXrVdV9+D/xz4dBg
+EPwEd5+IUlCkqF5HeF3KzU6iTWY2/z+1P88a+SYniKjln80BgesU+vmphB/2mJG8BRhsdp0Pho9
cnO4kpXDhGQE1wYC8iuF+THkvoDQ9M9mM2aTDSTMso/pIlQXKGquU0/a5DZUmFe8HfENxdGQb23P
FUY+o88EqHaqo9NdSuK8M/xg7z/hXTBbM9SE/hk16UCyYcy6KnlAup3IRXGwzyAAS4aKr76oAFED
vBGrr3pbXSmdYojhp9sra7mPcrKXdaRUPTvBJcXBUnS0VTIfp7WVazyAfRUk005gSx4ivwQnJnMY
KstTSJCHn4uf0/+zIsRA+w5+E/R/ksfVJF/ibrfn54t61OrpZ+EaT1PIC88OwhdXfkt43AlWIXEG
CoQuGf3d+txHGUAanp2Wai4Suorfcn6tRccVimQOiK5lOea56av9onGfgb+C5gkPIxKcTQElWH7I
JzIBLISesPWLVuRtMpHmeCK7jWSzKZ6J5BU6z1ZDzWiFGsK8OGCohbU+rnIXqIMFQVySrfGuvEfB
USsJT2nfEBGDgw1V518bxCtuCHVITUY4CL2pXyIptSponicDfrYciMFRK43W8ogy1VkJxlRobSmU
ISNKSoDmhxbhghnu4mp58OY79MM8MNeNOe9S8HEqnFScBpVWK4m8ch+VL6qa0XydNcvwWwGt6JOZ
uRLU6faJA9Q24yMtBmYYssGYNe1sj07F2lclw6O3kteFZ/2//1NJsWG2cumrJKDMZLPRKufm0PE/
OQA3BCZIZoglZLtppuUKD+IZRdrXXGjGmPTuKUeUCRLwAEq/l6XffAazD2+cxB/U7XXUqRlvdpvy
ufzSOa9gwenNkEdv3pSkD1qmgk6WVpZDxSs76kq1o+Qtr0aVeRp53P8DoOD73V0hkdpBB/Ylzne3
z332L5d/aLtr1M894PvNw+FU3JLhnsYTFxAnXuSCd67EVOx+9t2NSlyu3YEuQ+CbjGXN04at1uRt
AvGJJE/Ujy6Df7RBlDiKUdNgFc4yVUuLkURa8/+kQHvP/aXP4zRGQqqrymIEYEOV8v3pV7UPHfWJ
ysRleZp1GlDX/WFQSNmEAsUDd2XAaOIA/0pSi+v0p7B0ENYSjdpET1hR6MS/kg0t755n2/nhYqhe
BksAw2VFzYNWgkPDhHbmk8DPkLadVSSYM4rgNfqJNy8fkDoLt65buqeiw483h6qtVbE2MOmPJjn3
4uAyfOEKLuCQft+yEKo76fLFtB5zyPAvTzdx2tXbxwPub+swg7xAtWwXVQ6CgcjzEBzqJRvUlPER
i9LOE6ISJJTSJRqIM3dzACrpL+1FFjc3Vai1G1Y1udB4apm7CS4tE5t5rza/h0EBHppa0Vy13/z8
L20vj1HeSYYoa0OPfZhgg2abypWfEBcuYtI+9Pg/hDApZD7/5n0rVFi2TSU0tnagFmP2+sfWKyNs
uap4ceQQPzxqTq6BDOBFuZRiGprPGD7rmpCdnPIYTgkp7kNROdtZ+MMYqgCYFhb+z14plPoPxbX+
jdqD+3gjxMM7rYI0maOaMP4nt5ukr5TuyNs4Bubf4JlwDi7/1nWUQrBPKbQ54LWO1/I2ScGOmF+l
vwN42L83frE1MYJHgjoRBZHUemoTZkXCBUhyxwzd7lQT0inlNRra9ONxYv2Lv0lSFtcFUbR6BbWH
mjhhecL1kfq5CXjjcMRgSsjckTa8RBip0W1AzWzwaXBbWoS//rHxptAInTlQP75ldXzFuJPFmGAC
PPNKrJlo5bo8kvLxbnlc0lGyWMlV1gNGbf71O5OlHZuUVWV2IEryccD6jERpKqBBNjhpx82AQpjz
/lYRzjPiNx2GYtQrlSy8JF8+8P1KLECC+xMaR9uTKDbwEiogPcMgEUnl6rzvsjh5ySatgZCMs4Eb
Wo3Acrs8Ra7D4HoLC6Gry47U+jg+4XR4m5MJdWkl93jPaAzv0BfrTjhkafu6tcGT0juTqdxjmKA1
B9Y9qPvq5zBiGbY/359UX1VDNGhTSn2YRpzM4XUb+4ea0fOx3evvXJGsvBxmhsG9gdCCeT4wTGZf
Q/ksvIUvg2UqQX4t733Iw+TVYqVSq7toA9jISChLhRHSn/aO8Ai4PWS7kYTldTolPyF3mi2KoT5g
yt2B5PJwkYm7Rz1TcI5T5Fj6LXQwbR9lO1F6Q4wiaf70JRQ7yRKVoJGlqWD7wuE+JlLUC0LzRwBo
Gj2KEY1cCbPEs+I7zrq4Ydjrvq9fluyaYUoFsV91p3lG2JLP268yNmwO3hAKGPrvfnYgo9HalQ7z
DqNnSbPASYgtmSy+xas7AgsPCDSRS7TrqT1nPf4MTDABaqjk0QENWBxOY2MeW4OOpOaN+KjbR1gb
YhPr7DI3t4MRUKx8m7bs2xUQXvv7wTmOvCZjrGvIpgI+2uzvUGVvWYla1h8lChsT3Uzljt4IBRQB
6sSPeIRIKSWqM4Ud4iN8y/hGdWxAkJ3WqYOCWmS2Yy7t/qkHQ5btFA9D8sxSCUBdAH5a7vQmigNs
mKa0Hbq2y3CWXfdeyX51b8JYrot/dOB8Ys3epU4/FZwpJHN/LMkWVgfFowmv1v+DVPPJHHFQZPs3
owr6U09Jf9cNyUMDt6AQ9NfzuwaXHNjWC3FmqYh6v65MhQjoURcXPE//x6hmDDgmbdhAssQrCPkZ
dkd9WzmjUMOoq+y2BpBmMdMPnrz+i+Siuflv1F2GcZeaDnMCMH4lN5G6N8dJbtJe8AB7hZ4nP41N
N2qhUYkmNvDLxaggS1RpmTi4ASbul8xOLu/FigxNH2RPtRIg51bkrHXXFHq8NMHV/8N1tHMhkqMo
qaWPmAXz+Xlh388TOmR3gpGzA5xPMCOPwY1GSqFMOHbeoY/yp4e+Ybb5MYJNPOyOhDwY0lroY8Tz
hUsJr8ibBeIvLmZWLrp3gwA1g/lQM7NnEmA/7H2ZGBm0u8EquoNH6bKNe6BrVwmdiaY2DSegpzxo
fcQy8TrKc3AnVPUGekiEzQ5SOMYQAGU1vqiawmcWNshzKKqhiY8SknOi6nMt4om0Z1dhh3bclkW8
4SpcAN7VCkLxoPchfxOrFiRpxjDsFif0XY1Cycr6zS8sQbIvEEd+r/09sWoW14wD/B55ez2qHACH
U4KNQoN/86Otm3MBDW6GKC6+AvpHYkktPTx2+f+Te7+RH5AkjMMugO721kfeTagix92y0L+yYpsN
cM+H5RG/2xxkx4afR7rYLTt63hyH1Qr55s4PHJ8+JPh11RpUebSSlDGc3huDWeJCPS2gJ9yJdNrW
87ukV8pbJJsrTZs/A5LhSPro5IhzageF8y5wu9flAJPDbijaeP931vFpBz5+G/IptMakTR4wj7BJ
1FT7hf9G5+XNw0IrOdwQFdsDnBjIYPo/mtTsBb54Kha1g+7ZzLRg4dOc6XlTNtEXO7vcPzva1Ma1
O5Sdozpid+PJjFH24vTYCQP2ajMa357taQUfn/omAD1TVHwln3TgxcfUMLznzLwkaWCimgfyNrtC
KMpxxoHm1Np2bNYY8aByNx1ybozVjG7bLAJPy42UCW2p3UAyEUPKAac+Qmb3Scq2NmTgBR0wDm1n
8KBJXz1FwTR/xe+t+luIL/TTP/i9xYyuO6c6GyVTNs97ixWRCoYsp1dyM5UR/+cngK2nX48KbHUP
EUnyqibplH0KdYl34alRRo2QCKjKLtiDPnczOp68Pg/SOUDLqMY0sanKZcXmVbtXh/tCNEb+Dy6B
Q6Ck7NQYV8YTywpphvuK1wgNMUAJWfTYi5nHKRFiT9o9mhalSOQgOFoz87Vqp94MrIhyOfe9xJXW
gZBpngiZFEcGLSx4qHMahnsaufI4ZDKqxc6Hgk31CHv06m12MlumVOohLklzZMq3u0utB0SvEf/E
6nD7NfF8Vh0WAsLV37z0doLn5AuIh9RCFXqRKhJ1VMay9CUly0fUjlI41SglvkN0JG0egixt5Wch
W2wK1czjZ6MD19afLHMpOWCNNGjdV9r5y1jlyWNhLz1cEntLyc5CN1LULYuIDzyoGHex/Rj1c/37
qKO18ql8rTwW9Ax0nrRLE3rJZcvF5SdP4gSSR6sfyKDf/ckT7O/l9QgNDuELYy2mIdSn0cCj/fnW
zrIzrU6lCtXq597Ix9uBZ7aqa2hZCEktI7aP3oBt7G7EfROV8QBn3c1zBVYBnM/HoSIMQeyBvZlU
KmFr8iqxfiTsVj0GTtHjnlIPlZv06yw1eGN2YgAnbI6nncBCfz5s/PJK4f7KbES+2o5JfMQKN29b
40iZqEb6Q+ktkssisgaq74spqAuf179aFt481g4RpEjkzw33b+sqV4J3CmsWP7OW/QDkj7znn9M2
lE0KBWmk/idwLDPxYHW2wu89UoumWukwP7XZe20SWum7y8BEqmUOHv+i29GTluwUPnfcgKpajtLN
ADGYcrGZxqhOiuXQBAavO4K7vlra3T0hGCt2t059u+l5BT4JLWm5nxWaWQqlcjPlNi7muFhZANos
pbT6C/ji/VMAJPvb1pisx5rY++EVncCGxAwrAb0sY+uA3EtUKtFQXZVZ78t1lOhS1Q9jxoRHOnav
poIRQjsahlzxh9YbCw8nT91pcv3wAoA11IN5dKJhm57sFBGakSO/7FwXdU0u/+NcLcCWqJrViP3w
/NFMreUZyBlUofvNBt/cJFPl7JAhiFTtwFUoQpbkb+u0LR1KQQOIZcURhzGJaD0xxZULPPyRSpfW
8i35Cv3ZTkxVHP6QUQaBtCNLioIjS1REWVrTOW7IFVhFzqewWDuQJq1N3IKL16/hY55QmyY2q8vy
GunPJ4EJ5Ao3m+PrC+AqDuzygWe5QEhdpPYawxnU3G9T3ISGO8bYlGkQXOiRRmxFBdumyOvccePB
rdvGt5dDXNiJCtPNHqbNFfiO9/FQWQxl5ImMoRGEn8ihU0v1Q7dwNLiWZiRkpmbL4P9X/kRcGMhA
1mxCItd1wtOmTkv6OjXctY8gIx9O3fBK2OzmYPp01JZ4OCYc1FPhedcyVv8NPfOV+mk/lVStUvRn
HvgihjXMvS6LbWiXHRuRmlCWv6n2xfGIzvNSEVR1aJJhwTSV6riBzpqcenOmneEO3GxgiO144PiZ
iV6xJy8lwIDAFhzMMfaGpC8BOoEBpYABDooQBDVSySsrotZXKsSUtxv3j/+Wk5Fr6g3mNZeJR8Zv
46UBjA0BIsl6VPAIAYR4i7qqLD4e2Hda5dTx2/nlFbETeeFohK3yW9KzlFCW7Z6L0/YS9GN7KnZV
YmWwjjUmRnc4XjWK+XRUM9kfg6e6mEPEJfCY54+X/4NmWVBAeMjm58tv7OCmk13JHOTo4TIB1k+d
OyxsSPIPqEUCMWWsimPoEtb+OH4ZX02qP+wTFibqLbs9SAYUUeOnUj26LGKhU1uzUF+JrSQ/8D5C
kN9+0rb9ssUmz1swlngff3dAmcO1pNeu2+7je6IwfGVbI+lI/BnFghbcDfQo7WsCRZygEYkVwAUL
VtXs4cLArVQB5aCu/xh+ZcflGBaD3Lq778VNuJT4dOljQM3eClNcCX1vTHH2z+2ffp4IBR2gLGn9
aiepxVxyXPAarqfOD67+/sSBK4YBbKLGcIM7hwUkL9hsIgcl7HEtQHZYp1N5xdtvwQReNTlC3OSu
lld0TBMWPqt6O6FrRLwzk3i70aztfE/yCrv/P18Yu0QL48XgqSkCnak8BBu2m3jZBKnWKlo6LEMp
uAiRAKpN6ATxjyR+d18NG75Xh/YAwDjFsRqadbUbR3FeSoqzpSbYKwMTP67NLk190prRqUtPGULI
Ve0zRZXwculqnfSeenlDNr/lR8tGEp7MG/bZL9oWl/yUfhgrJW3Ma7XbKapJOEUDYVAfyDcRgKqQ
C5zA+L9LGisb0s7473a8YHaE2r5R/BnZo79g/qcKtitOTzxm/nKVhTAMxq4/5FbbMoPridA0TUZB
jxSFO3OdDuqG2ImRSAApnzTUvT83z1outbfQImRXHZH34JEejrcBFCg9NSsKHLz8vDBBhi1NANDB
KkcBxOrFKG+JDOEjEAHpNj9iO2G0eGHm418QgXS/G5tWOlSfgGPvLkxTTf7N/tLNGUMJxMZx3jW3
sqQV/O6TW0s9PNKOS28yINbre5IYjOMJUOJCWXLDOkpIDaEiVC4kHyrjuIu6Qc22pASR6JBy4CC2
dFhC3RrIyi6Jeu5TXHuutW6Zme4fLBJfB6aLf4tj0LYETFtbHzk7SwLBsTzdZPhXmkWXepxy95yN
a3oPUVjQGsDSsqhcBrLvkNfR7NZp9PBz23zkNjZvXeNNIMIioC0m0L3Vu4trTSAhIL05ewnxsM08
3zTG9ai9vFqp6MmrnoyoHRS5CoDE4r9jQsUE9rD9GupfV4dUf+DWm1XmoMuv6N9a+a1LrueV7eno
sRP4OIilef5nR70nCYehgq9drT8cK03HAprVN0K3jgs3jJN7TEJoCXwRxlF3fpIuECkUCUvYTgZ7
NcjGw5DhjTIoigxAW9duh3goOWD22NtS4nDOuA9K26ZAFuR5O6vwKMIn+gzENlARFoZ3rLoujwlD
H0Sf1Fa81YcDf8B8bnvycpuOSi8JF0P/PB9n12mqa5mnENVvJrfYwGTTN6jVOnYN84SoCv12gcTi
uDkxMRp+kUqJ06ojUTddp8To8MAnkeyw3AZ4TAWM0iVG43ksNyxN4Jau0wITq/uIdcVwaq6zi74C
WC/Nb8XD9GZCyqGLpm1i/IkuZ5vTGoZf444EC4Hh6x8rAHRkvY8jILG9/zsw3RH5etn3pyehgYmn
DL3FX9W6wfGzmS96doXcWokSIsK4mPdQK1n7rojr9PgsO6Ij6hKW+CdkVhqsJi1jFdEmR5JFoZxP
1Xp22ZzAbs4HCamQCoXtqC8055Aku+ZvyJB5DMlIQIm2BJ3Wu7vPHSX9idcTaSuBguAGVgz1fnXY
bwtq1y80JJO0OXeS+9nI0MkYZOKXGcGYIRPBx6xC1+sVDgToNxF8iWD9h9n0nbZ4V1zr/ZmLbkvz
ahDMJVDs28GHQs5cRDYkjwUT9UxtbzZs0n9QUnb4bjUgcyLP3ExLcUFvujmqP/oMgPqxqp463PXA
e/qOcp56PH1Gi6PSwxnsgGuqUJBX2QnyD4ZjGQnfJNsIlX220qCNPEKrt12c904Zbp6c0M6EtM3F
W2ycujqxKf3fbpjXOUadx14KQpReB/ZHBX4CXkW9PkdJCzrC2u+Il5SNhFwXvFEKZlIhP/NmbDRI
uHrhsGplo+2OA/K4zq9jDZWCYcI4irxk0iFM1xnSI39qCk9hfDfdpETE4i0Y2wl72U+Wat7NWfnW
X9wktZvhZ46VQyKYne17ITj6sKzSEFMS2IYZAbAU2eRP+dlARBlR+QnBBgyEExi8W4D5Qlr3ngtd
2o2NiIg41P9MlaBjT6YRvoDiI2Hjo0WpUio8b4noRatSpfTbmMiIBZE5SKhQyGtQpq41M7WDPTRB
6E/jml7ZTHjtqCmSh1tC5vYwSSw2EZSNkHx8taSm951Q49zOcPMErscIahuAVUW+uvIir/heGrtH
WVz5Fjp/xnBCCzD3F/nVYqHQvimtSAR8pZbgwnLGIgtID2RTDqlk+bDzKogNdLp5hUf+F4iK4qvf
lqxp0l9S98f6UvCFgBd1pyWlUF/iIpzvgQbLchWt20GYJ/GSlPdwj57SFmMBrgCd79zcevqCd9MR
DGutsajFvhbk686MnWAalvyi6AgO7XKd136jbyGecXxiE7UVoybw3aP1pb4D0tELeJ2zT1jtQX+u
cMHb8Rvds5Tpo8zyaiywLfg5hFVFWWnwbeOnSOVBEtQr6ssFWCuWP+vDTNy9Zi+x5T57Sun/SWT6
ZVWcLT+/tur7uttb/AJtGMGZUkLy7aU/ORu8Oeewzk/KgKN40aYD9Gv+xUsuMAv1m9/av8R+NqIo
c2gh/d2J5kq9R+oJ9RN8k607ENx9nEQ4MVH6uICIYPElkKbtNDrzrqk64fz10I3uFmUPWE9W3owJ
C8Pt76ZG0Wc0w0cKWqep5L8kI+tdYqSM1akxOpkyI+yIGXyU1N1k8WAgwJvw3DM2ic+ERrOdmZmM
Y0xWLyyeLLPBT86OIigb7Q4pX3SrqM2SaXgGtvzkIipPT8DKD8mgmQDTumtE5d8afv6G4XpHa5ZC
a2mvAsGbkmZt0QwEvQoCY/zpfXOnelM9Vx0yK/OfX+AiqU+D5IZJcDZIzDlwTBWWcRFGHaFdYNNm
DilNi3DlDq6clpJEfsnBbpH6W4sm4Za9nXbpPNfFpL1w0TKSiPmtoH1CBqGReWKuFjRRCPjol4br
R7t3Y39+8JkM4eg+ElhRcKxGi1KSwZDnfIFXwO77ev6JQa8o4QDXDECsfmg3mxVEIS2JqRlXWeOj
lCoVdyLsXleoKEFUmCaeYYKSKzP6oI3TKQbpUn4qz0woMrmcPcoDqrPQ/NKsQE9Q/CEaln2VqmoQ
qG+d9hNhAwhZVw/qeIqekSmlCXwHwRxgdB42vh66/Q96F0zP+KpQhbmss2zIUeIKW7LN6lvJPBs5
7xqdgUTi+GVWFfHFEtKwGy2kIy99d9iNtwyl2NEMs9VUGcljANsswGHNOd3nZbQflcTlQ+t+/t0g
dnTX7uKxS3FL8k5A2A1FAiMQ+LGvIS3xLrjkj5jDWa1/6uFKKoOkWQpa6eZBq64bivw1nxoQBflp
LIZrML3nnPNuiG05ChCUXLiI0f31LwQBWBSMjDyb3A65M+bfOD7HHUNL4+idzT6MNYKmYM1IR5jC
RY6a2pCosfOmpeGfEK5XFSSRJ3auDAwanzdBiA9H2ZL2EyXTMVWO9iupFWqMbjbr0w/eY+tIk+oP
s643/zo4UXWWgfoZY0Sdnj/gO59EjK5qTX7xE4MldlLuog4i4HVwau6aYEUGKAwrNVyGbLAwDl2C
SxfLym8j9mas/MpTWvphrTEnspZGjLONG5mV9hM5lMMihyxYJnb8c0cZX8EBTniyQS+6bbckEK3D
rgqdxdMn34JLxcQspGNGSsLrs2qXt9APIOrZsiGSHyR+j6h2eYYuYgu/eaZj5aIzpiqe7NkRoSxl
i+8bCUW456aXXk2WN0VO5ErQLs0eDtMmfNAt0PDvMZMIILw78m95+jCUEUCmKLOXSrKxkaEuz2+n
4Q/7V1wxAk4s50sKn5hIKah0d+5UX9GXROA+l79FlcwWAEi07t9RUETn+PoAfrAgx/TaptPUsVbG
yHXko/IBbjP/H2H/qipTBjnloZBpmbZXYwd7DAAa8dzTUdt6zrbXYGlJd3C+VWODxqWjpDtgV036
bkX5XvkFq+EnGfzTEZ1xmztcdwJfJgrVp9Mf9i+QUi1EJrnhW01MSvTjGaGkjmrmOjTE957qWZrt
HdLkG76qw1ah5xO5P9phi0i1pdyfqbKZDqvMRT9JvWEse+hwdjJbh3zicW+3Cm82d5uCbwUd0Cz2
TVmW+KD4jPSe+iv9SG8yFJngQrnVz+f7ghdKEHXqit2Kg4+nILYUAmHwCkZXpfDlAgVD60TEIay7
UlGwNq6VTTZO5rHqFLnT58sloDlQg8J3JgdTCHUQE13z+6CZnnbKQTUcoh/8d1aN6OE3Fidq/vsq
ecLdel7J1UgE/A5Y7bFVVuWDdaDXFpCDODLuqYk2rhMONSgCJz2b5slHDlu1VeHDHyZuow7+4RsI
NGIpO48p9HmqmAjx3Jwf7d4eBq1kocxvQXZZqacgZmniAbAEPLWaHvRPf7fMfoYwPJw1jEOrCo3H
z1q1aGzTpepgUPqbjirUvs292uwab4uOPsQoYUFJPjTmqjWZ82f++QmjP1+k2w9jBtwfPLHkwyHi
1H1cXWVGTUNy2/LpQOB3L8KTfRYPH3tvPJumuYXQQa1m7UmgWGJ6/utisprCAE6nUzyCpna4th6+
X1Ojolmsy3P0B58BKFSF7oNqaScKPKQ82w60aJ9+GekH9oLifMBrkl2KH6XKhM2zNb6ODLd2vTOq
a4bhGjpyFPRVfvl7f+vsG80cyVxH/efWou1nIRDtibd+TuWrcT7ECQQtJg8T0Qd/rQuZ7nvJvtX/
IS0Ktw62nCDrPvhss2OAXxnJiSxLZ85YIUxuAVMRkkyR02FQtGN9TJVxuqojt/w06DWRIr0LGJtv
tDEeUFKe1ZuRpDFoPC3TDwnpm+tQvYCkZN7uL1tiFQqOWa0OpbCiT/nqmusw68MlE3iCGXWK5iOQ
Sh9hcm4yiAPuZcV1urv2Bp14gjygApBama/Vgeds6KOGOU0c2K4tbuA/N938/DbxEZsTYsPwKBQn
5+NGnSGHkLncndN6WgZXy63ItDeJjW98OZIkrNmFzEzg7CEPLIgp18V7cd5/+b+In11UFjKXu2WU
zgQPnWTeNYdKn7xBhd4SFMH+TRFH3u/nJoWi8bTSHkIh1jrC/GMZUKG2lSa3e3R8WBOHyXJHpDUY
N98Zw7xdXKBTTNhxqyH8oS9WmTK2iaCY2qyUWREhtlZsAgfBUqw9DOEGmh1zHCxIrjDgm4pnOgN4
gTXvczmd3xzUOF34h2RYDJb0YIFTCXH4euU7SUXtuHYhPxXrTleaL5Kd33bogfYu25ZUZd8BOxQ5
bVhVfQJ6jfxtPOW6zjAFHh871DTlxpC6ibhAEVADNYha86NE5vNv2fy9icvghWDia/jxLApiISjX
LLTbn41gaVryuLSveDMXYysJXNtLfvnOnATop+N1C6ji5kd8zUtRkX24hLdBVk3rNu44dNF9d66O
FHe7qAKK0eC/QIIhKSiY0nwZPgdGbjKhYtVPgAUKc2zMMuvp7Bu9FLmSASrkkrhga02O6182sdIP
5F5OELi836XbFYjNvjzbO3pHTroHK/aEw99PgiPpoq1wRZPwbNzGYxgSvfmdPwlmsh4YauPcC/5v
w0kXAdJ1g2+4VaQsVtir/5kLj4UhMePIhZ71BpcED4si9rdn/oEb+12sUt7bThs15hJH3Tda0tl5
WYGohN4sU1Rdu62hzozGkPLOnLl5Dz0FEafQ9gb3N84Ik+W6FjSodFRNnEOWwLzHdtQW0oCuGHO3
/gZ9f/pmN9Z/aP3q9gDGl0dFnazaHh/oyyN0ZSNpUScuoWwTQehYdctJWqmkc7VWa+WuOEpN83Px
1rdgO6NxAr4Qkal6fd0eOf3EPBOcwSo9d4N3V7xMcIH3SZMtiC0KpvVGLtyx4yZc59bogmznYLyd
pUxISHd6tOmAg3nTqwTuyj8Jyq1DUraQO2oJVHjDHPUhADcbnLuwahtX90y+jm/oNz/jb8wFG38q
R1K5HD+3dGW+CqEvvnILcn/Brtt1h8N8GDPnfhfQ0XSkfOvB8n+W1fuZqV/cQ8pfLRGw75Gvt/md
qAUS3zgIsuPZv2/ZK4XfmVJZ8jSPnXEq3FCYilT6VH8Ih1q42TvLZ72r0Ap6jTf4kQNRbRiY3RF3
s1/MV5T3iXM10HOKjuZuSW5g3ZCp3lAJBomigp2RzIK3rWyO3LkdUhalE89H6ogVQaHLZ/aAH+XJ
rzLbey4WoNQmq95DaeyHwwbc4jlRm0kSoVhzpUdU40oQ6/+bxY1WiFjM5a7LSNGMfIBbiZI34vLR
TWcLLJmneMzObzB5GoJx14piQ5C1zCZ3N++LIRv0JYesZR+8Jc+t89ZslKEOyI0HPmmcAntEpT8l
ZPQoTkNa6K6BSoX/er8Ff3Gcp2MMs0gbKZbBWNsxrGXfg42drXWYDimC2QlawUwaHOe6c+D/7Ql+
4jW2VFtLgYOpThuEklHxJuekiVSZ+e+h87d2OFgqnAXc9fVpFt6jpQF1JDi34bsOIkR4eFdEIaJO
MMuIbdzTtHVVMwmj4FWJHOhP9y6XY2XM359gp2tLEljaborpUmJ9BvVq1cmqkhqbNtVOS1AD4N+G
lF+DtKN37RnTeSn4Tos8BYl2aZlDtFoxOgho3SZNfIXUvLBnsZBfzJgoxuDxk7gYupxhSm45DpfC
J8GbZQfGDrxj8XPEkhm+PPDlWo09gWap8kBj22tSa02xnG+cLw1zhHY5rKEoE5tS35sfkN8V2tu3
HjRJyd/R7/56pX9X7WJcwc+tQmILdNxRwlh3mhimlFrJdek8vXFqzxC3in9Oa1vpwRkTynhVkw5c
32ahQF+8k0WM6LEmi6u38ySyN93JdkYcaWlnU2DyuHZd/D7G3XTRahpq3nFJKfspasVx7guj351/
sfMP2+XpCgZ2PCONi3pv6AQ+ySb1pW3dtIvnrNlUGkLLfDX5sTRxRoyyhxlVcYY8z85BqZ6mCG8F
NMpOWmp2Mxr/ESjBoyOnStlJNVf31hmLbKmrUW6Pf4vc11aW1LJery2U1SkrQrZECZO6M1rJlIYv
uC+Vcs7NavdpbG1bC3fT1VE4xQHCY7kK28YiahXPIasrk8qvgz4ouAJ/JHMAngzQQK4He0Dbnu7G
8rvyKfDJikxgaz2Ej17dv3dCUozzz7QW3BTaN+9/e1ih1TSspisOHiSFfFWeGnGNlKgfvGz32ixB
J4qEv/9P5wfO52hcvEBsqABSZUjjW7ia/6sVWNzfYK9utXg1iP1Oy+eJNWMytCp2d3RnOoZpCdCY
rM8DLQVL+LHdDB1ce6pncr4RoGq1hoiQDNUqx4s4LW8o2AEgbnoBMI9fFZKMkgnP0Whv2A2XXguI
vNM62woHQkjDYsbKUcwB4Dyw48Ch+efia8Fp/HZIgDlVWws5OaDqH3pM+d3bb0VrTn0Awpwi8uX+
VgK34zgBdGI5mvUktI3iGAjdkrR/ua0jJmXHDDJ3+e5BCNiYRxP5Jpk87vzGco/Up0tFJpegY7tq
kJ1TGAlxl+4HBFRaq4QU+dZjm8mURZraIIsDbAqCiRqju2Sq9oQImSiGq7w0zIz+fC/VLSQwdL5F
aftYEVWt/1gcZ8lzPdqv7AstMrTwzXDzrDeZj4J5bvltVahvhSqQxJBK6fTy7L+2prDAU6nlrKL/
jvTN/fNm+bKfAyuabismXxjODdLdBCDODkW0mNoezmMBk6CGpvhB/fxODORozdXWBXVjtNcnQsJ0
kI4EPrb+6oNfpfP+ggzvISTEGaOWznejrp/T+4o26ZWSvZ9wrtUKrrOGrbPzAmyHpGB5IPFD8cCO
VZpReSVN3odqhVzAx4I0okfkkpLgr15dyzHFvjgiUJy8LKg0odIXIhM3X28U35gbPQSGJE4kiUhK
eTRq7h15Y7n4FovCrRXO/SOI5pw86ag84RFJKevI3yBzlqvn0sZLRkNDQ/QxUZ25QS04A6l+kW+u
Y30bpJAySZ07kkl2M4qH34OQ5pCQRt3KDX2dKydFVia6hDHTJY97wpQTL3ZnDKPRemFTr07P/1yG
7fEdmVezJfhazIoqn9me4hTJKVUtJPP6hGyOWSAKQsRlWF0djsZrpp6OH8LaMWVYfwd8+kR+dfd9
sfyGK518O4gzc5tBf0CZAjAsFFiNSn37SAnNtIVVZ989qlLOszjNqnnTbgselHPEbw0GU075M58F
+OqpAgRnLBk07CC8bbeUSv0YoV49dtgGgMmMhASSaStsFiO3wro2g6tDVt8E9Joh/DDj8Er+2NU5
8AEF1TFbyZBx/NQ5OJPIo4uO5dNLlKbyBrPL4EOqxbkDCQOpiYMaKwidzl8rEgox0YY5aSozXm0n
kqPq3YYDMnfgncq2UcRXiy+iIY9D7yyWZcLrFOwFQcgKSEt+z9fba9Sj9nBwl8EEU8tJehcOXuz5
iLxcqsIOYEIZ+azvr1QcYtsLlJu0cvy8cWvPQkKSJC7qBIGgxXOWzti7X4+1bdlM1R39ym3A5FiJ
QyCDjNICohLaXbBaaTLHoOKd/72nRNPgG4lacMflW0jbuR+KumeqYFrc3lRmKLk+Ozh92enl99ns
91A/m68iIWs5CQ2GeOTdfRILvDCCYHfVSHpsLs2B6CXVfim9q4Fls8dJWdOEmmhjfhm1xbKr8A3A
8Xu6YrxokPhkGs3v0lVausqJuP84sr0ic962RIGwOXpPAhruYf40JfgOil4m5/GjHe/cNQwAIJzm
dNi4ndyLyeqhVYNB6p3AbAqaVd2d4EI1tDFp58BXADXkqD2dYk152EKi0rUB8HERbW2xW6tkP8U+
qgsNFWpmP+dFJnL7eNYa7W5EElAlmAXgnGbKx0hgwBVvNFRikpYxqVAlTWdYJ4gy5bvXrlFBnuhH
i1ojVBoB1v3xRGWMzS730BTFTWYV7gAos8Wt6R3jxwE6aPD/QumCtno0HgS2M9zFlQYAl7jSjgbu
jeet29w/scXLN4gN3af5Vske24ZP5IQsOZGsw08QKgVY6OM5JQK2YBAzU9wqL6DQYhVeHLk2l6Za
HkcbHyEaGJOT4QBaKvLjtj52/fIWVvvfsMkoQLFr+LTH4lATiPatHstIEmb4bVDhWg15ot1ndd25
2blZmiZk8KVFZwMeXxYsXE7uOTvYEOkPKEkcbU+We0YYZ0JXS1V8lbmOUVM3hGMI0Kv/Qw6s54ka
aN3UyjcbB3jTSW//KB3/XWs4XEknVLhNAju3DNk7lOXpn7t6Vd+o6RDcs7UFx0/9KjlOzkumYy2b
7gmKIPeSB/2+yicwfbsBylfDEmEj2sS8ryMQrYkOGDwLgYZS+wHp3/OytIzMccoX3XhfeRrfAF5P
hoKCSR/PHiW6UC2bBL/GSc29YR22O6O4Wt2Ro1tdNNtQEOmdoIuT+YgM0rG8AxkxGUylEWTOb5I0
8AcvBeq4fG3cfxRrcEniOIj6pSH5RXu4NIb3YAjaLagngWtKNjeHjtnCrd+oucghP4Uxha1bg65l
1M/JetJWvlAPc6ShXitrzH7pxJoFZSzOLtepx5r80+gMTHFABmIxrhFnfdSYjkvXbqG+oPZGveit
HnjYJ8c3y0M/MNMlhL5BGOxaJpQk8DpeUPQtAtnb/9Sj3WwFlf7eZo45xV99ebp9cUrcLehCuv3n
O1PXLTlMkE216oc1KNuEcElx7tzPMCNlvPF/vNiHo5ZsfOFIwM1eJOoy28GjRpUUuNl6JxH6Dl8+
4zOhRWiosx8UiAYlN77dvHkXXNfxN5WOglwJWoY6++OW+mRgW8COzjOg974lXs262ZdaFeCsOUfP
jIzuZg8IyftdtzEIUIR+cDipI4P0/XQsB11cz/1TtIp9RgBKs/bu/vTIlTWjvZFRhEjQi2riIecJ
QoZfExjnvbvYyOUflnXmweOyA36IFKgoORUQgwBKwOVST2E2srNVGjEMpAtwJ+zNzDgE7aujAbTY
1coJjh7sWRi3FI81ctEjFq1GSI3XDyUgJ9K3R7stbpQW/jJgGy4KKXOtg8SW1agT7CbUOB1e2PJU
cVn8oDtzAiI+KYcNDjrbldM3ZSHI0pA4QVQxEjY+N3zARHH1/DDHLNQhB63To5z5uBLfRrk9tJ2D
NVnRcr0zJcT4LYlDcThPO1mjDmKN9bD431qF7+U6vNjgxdzNWPV/6rOz4/4Osq0CkkGC+F7w+0/D
Ou0YvYZXvmT+qIIg6/GO3IqweJIIikHRUkdHWLfvTSLl5vEfxvNLNnyw7XCHjk6HOIewdaydaxds
dEc+NErO0bqTy/5cWEwmzvLuS5m3bJFDEiA5IBMlVsJ3fQGMuDrqAqzE+uObYjnbXh8Gz9nQCWw4
bEenIeTNMkt6z0DzyqspqWvnnzI+U31CD0TeDISNExWY1vrEUr9FNJQO22kBTpxyS2TjOIM+kWy7
yF7V537fYq0WqAC1DdRxdxWrYYEU0wye22fDD/gOj/Dr5Qsa/Te/Ulv2YoIM/YZbvF7C6KBgY58X
Cb8lgLsHG/F+VH+yXrlJpyi6+5v+CjB1G6Qys5IEMAcHbkGpZHAF6EE15g33SGMSxKhWDczmYV9W
L64aIN8K9a5vpBV8LuN5r1dxZEbEj2lPs3qf5GU52FJDA+YQtFaRYfFndz80lsbETiJYNjlSwaeE
zVbSv0C1Ttn97qrok7FAJU8++Z9Rhx7Q4m/22Lavvmj2WUVgurVCTs54RMyhfs/9UWfFqXc8dguG
DV49KOp5dkrvU+pjCkV6K4gEjiQNdiHnUQMO/Us+fIWFJFkM1luFI2Go7qDre9yJ1jFHECCeZUso
d90qJAT6o1oCyXPqmK8REZ35b/Yx7OTKv6A9xgGXDWx8ldc6lkp/+R3LE/JVGgULvMf/0ZlSuK3r
hdP3qbnu+t/I8bkKzESlVlyleMYulLMn2XrSX+y/oy+EOZcCN/yd2AQFET2RX7SIFudrt44/Kdkf
/VxsUBRJUSVKUrdBOeTs7MHg/DasvgJARLldIDQyxNmvLyTE7hmoK0fWZCcq2HyLqkoTzt/t27VV
OWVZc0ZiGiWG9cXvL68Oi44ImTsnwhJqyS94ReVSNnU6jVBt0FUjPbPgyhTTh5LxTpj3SeA+YVOt
qt/Gb7dY4yJLr4cUzjYOc++eRagOXT3juWwM6cHn4zfUNcFf2FQUBxLOzucWRpU2nkZxzm5i8BOX
M45deWlemONd5gJPL3k4rcSgBX2J8J9HJ0dsOLRzY2Bjl11OYHJ+tfXcNyTgUjZb87yTaROx5Akk
C+JT0iGXjkCbVuYgv8sdXw0QuTILPCH9U/APQxN/dgjdm5xn4zXVC4I1E4RpL8ReA4XBHh/26xvw
nXbZkr2Mqy8QCGUEO+0xVX5AK6IAW3e2Q7q1SIJge/IwFjcEy1y2H9o4u6FgkFlAIp99eIg3kyaL
0trkTBbumFO2eh4YUHRG9a1z5Ld2SmYbs3xKR/inbnKLeCFNrOKXH3lqE7NBM8rRE9Oue92WwBmb
n01C50PYKkfFvlcrwvpPBva/3hSZsjkAa1azc5PauwnVI50DL9X23GWMD5Td26ug+J2XzI/Ge3Y1
cB2m+qT2c0gR+cpb1wX5vrV2ywbWbIOnMxcnWZTcwNgphNVSiQi55bEPeW9jfXIHjT2i/MPjDOMj
cCPmAuLTPUMLSkdGhqRGP4WeCnNwZVYt2uN8tiMwYcoYZrdDmEyQX3bO963tNThvIddaqEXKi5UF
t4ZvBYdoqlnoB6SKH5NuyNizej28ZGUXWOkg1As0BIAtxVOyWDNP1iVTqocSCyHVO7KrxZmgUWqi
f9dQ0jzU0yBz37Onws5RcWwRPN0Ox4PGGHPEZ5mygFvi+Oh6qGt+cH/tbjwvv44VhsG5si/7+hYD
AQv537fbtOcYULFjzLeFsnSHnf7jjYfPQ2VxYrRbGtNu9v+iK2N8SYG+E7q4rsyA0VIjZuajekdB
0Xrjc11QToeN4SZu8RIpLtaeLRVF7QLU/FeN+Hma0j2wBR0ScFFWKTMO4tRAwBxPISWc+8tNDlts
DdQX34TO1zbw1nIGoivTLlZB79NsoFdyFqr22L54kR4EXMhPHGBo9gIZe3qX5GnV780UmKsxzFn1
KxvrIylNjsnfIKhIFRPAUKQwLen8L2IvAe7CJ+o8W8zr6BIC7sJoplgiemnbKfCorUo7mRa9wTc6
atAXdpIKAUmBQF6s/JW7mR3eoXavGXZIls+key+txjy/Pk+jurBA71Cr+m3cDEseBAh0s4xeMN5B
59Q72VWcyDbQBdYHk33SU8i5uqVa985nrv0/e6bgV39U0OoEWZsxtlvvZKit9ojd57zqPx/EY6AU
lyIV2s+dZAeyoPRDaO+tAKQ/AaYpBsYvNYufmHlrg2Q6yT1cARQQJQqnOjNrsd4FygvD3/KV4xzh
OENrTYh+I69xo8qFWjPf4NijEPaQdiwttPQrc96UVOOQ5pnh0GVYYk2CRGRXfWI6nyiA9AvYMIb5
e3mrAqjWP7RK982/fyxB4L9NOGjJLjeLtek/PxgNgwov1ZQyKUkHBnz2GYN6T6fwoCYidLNu0PlN
lhBa3q9dQ9WXbi7m5xJu/1WbKu5kvm53rRnnT+tlWMlkX9heuJv9hxKKxfpj6+lb2Z20t9DyWv5n
8HRESzLg7kjAz8VA21vXVcoktfq8FVASbYR1ObkH+jvAGb9x3KaUqF/cRxqw9JyeGOotKImrmsyr
0T74XiWEbyoHO6eN7bqbtbQ9MxYdnUCTcbdhbaEFrdfzSqYLMV0o+XwKJh4o2b7njx+oboUqFkxi
DTfv+kXhw8KvqRAE7g0xLLDHu/YT9Ds9o+rz16ljtW3HwoZXJH5jjrBGHin5DGYqh2p7s64dHzq1
grZRmC6O9IwlMTGjzeXvCgOhkaXT+31pms1CmLc2PhEH8pSbnjnV5sJToO3vmxB5yPN99l2Cy0N7
7NzKPcPwuNTZR7JufUG0Tam0q/cA7DzGWciExu41JAOuz3qnLEI13gKy9wfacIz3sVAWS68F8T+Z
/kh5DjswAN7q2Q9+ZETyitNV91pUzAb6dwXG4mEbB3lZwcryTMEibmscN5XuS06QoaLC1Yqoq9/n
0yzkr1lWw0QhCIiy//d2CaIDgyfIKfCmSldLdFOlar8gr0p+SJFw82q/DY88AkrkKyizfoEHdXTx
TKGrPt3nceSP9t0BAhmYSFo7MAF7W03QWBrROB0q8VRAoOK7bEOtUefX0sJBbpKb1ek8bTPkjSiW
gLl7ZHMJLLs+TbC+LXjZfKQX6EWI8Fjx8kLQLtfZq22GwSkHrWjZ/uqTZEN9AoMyKYj3eTFjnTfj
ewQ+uaJdW8IfILM9khmhnn/ItAVk9PvisdDg6fB6MWhclsqsf96FpAqpsNmFYzhPSzHltkHXWXSF
l7ZJXfNNPFb1SV1x/Tn9VfLeclHSTXDNliyf0DAyScjly+H8FLmPgej/8kD+nDmHXJ47WjyzuQk2
yj/3APthNV/vSHtMGHyEdl7NsUUfB9WO07PyhhmrYD11CylWWoPjlBR9EskFqDVv/PWR5OkQgpTT
ZOy2G1+lWAmfoa/BoYFjphz5q195iLwB5YE/hVJrGuRc1MN7QdJYZjUwm7crrM1L/RTUeJ2yEjkZ
DFiWkkvpbiy5qyJlRuz0/hIyD/S3PMiJ7DJl5jrVGVkLpykGIvH7c4ETbX37U9AjgfKIweiumvZS
vT6aLh/tV9F6Kd8enWNsPcdVS0BvE2I4sF3tJZnE4FIJP6zVtzhuNdrLmuvU1IKB0xJjJXjKKDsU
13FjZ7p0hh/g7gUXHWthchS243AQaCiOsi1GEC26iAw8Ccm/9I23b/2/OSEWmDQcQE24Li4iqB54
pTV2EqW4DFxZRR5gaq/JbO6w5qDWZASHcsWU7JqPS5igGn1LI7oaIFMoDuXm3vuK7DqBbYelbzUX
OELUKjyV6GCwYoq97nYNQnULQH4fig6EzluIjyNKWGgc8dGxU/4u4zd3yC5Q4fArs2FPYrUg1oIv
aNXSsbigoSNmild44Cxtk+V6GmDz1C78mYubcZjlYGP3BD4aGpboYypbOMKYode0+3OPquRBc12P
jY0uVbkOyclRYVoTSdO4+HeXZklyhyX/lldCHMiXFrMFChylDS1AOVOzoQYYZ0G/UQ9wUEmUQCn6
T3UafdF91ErXv2RBXnq+Cx4mTtybF8jNGBVo1u0OdfCbHrA5ljEGkxkGZ6SPaNLZO0qYFzlTTMl1
Q2Yln9bXat8L94uOXtStZLULOwpLckS3SXWjaodzaje4pNDhbT3u6ZgKpxE4TVtmLUo650a2ITqV
Dg+8bZfcCHj2pw5Ku65OO/SsjERBUi8Ih0Qiuf0j88jPdGCQQw6CzfyMGe6T5i6+QjD54qubYwU1
XlK6rVAJ+3r1ndjQiAG9xjhw8FzuBopmsN3XkSKQPZPnr1lGPLkQnA6xrrWuzt/R3iRXluP51qi9
0W+RQEwFSzCrIFZtfoIzsOto9Lafmi2gg8CkMC6q+riKlhCD7TpkE3yXBS+p18IMg5+KTdFOQtc+
Lrt1yOa4/pCQB57Y+9feKMzOrbSEO5Qo9lad9Nc3yCGebyIXuhTm8/iqxNiYCQHWTFlk9G6fEkzf
ETMWwFo+AJoX6MSmcO5OlqGWrUXR9P76rtOCpVTft9ip/qTlMiPCQw6JE/r5cv0Vez9+JtmltUIG
35uGXOqodQ3J+y6jC173gyYPu/1vLPi5z8HdtcGRldR8fGz+Z0Yq/0b6/Bpn1ogVDRe5OXFZQYZo
VUWIQc0nwKlC+fa59sNlnC6Yy8x6Pl5rtRH3rrX4dsMc5Cg48UwYRjtihDoaDJkQmP/Qu3qYmHGj
swt4J1pocrchFwpvEWIvswI3LdAGkqhhSWz6ei080aggFkeDSz5yrhJAP65aU8lJMD2IA5DndaJr
iL+JfS0MmtWiHfsD33DITbaadYzq9+u2KJzxd4+r+9R5MvNz17jy5qROWcJR4YfwJopUORMx85M7
CL143SgXx4yBnuUt+ekBaz1e+fAKnFqPK6K3MxNLI1BC/quzTukUV11rFI4YC/Ct4xTYNflOd4u8
hUKIpUezckgiQrQCTrUm7aVPkNuzWbJrMwamDUVj5qdvMjDBeQDG31e4vzcEOC4yXtvVBUpyGqT5
bk7UlyMabWRKzu1zrL4oAmEhGJ0wJfCbOyTtOuHK9gb0xcaaApsIxdjgBZxev2rBfisr9cePnJ4N
Nxx1VHRO3qtr013HqA+wGfKSSpaVnQ0aJUZr8eiHqsS5PLVVxI+Cd+x6y5tiUPzM9lJZLrtSCfQS
yBbZJ8a+JA//kFPveNu3vVHsc4R/HH5KoYPlo/hZ7Fujzz5GOOwHckTXHFcYHKgFP0AmGC8cGQau
xEjpFnbtWD7lti+kDvFybjrGTiGw4/JaPA7ZoCz0dybSzMR/WdRl7c8YlVBWJFVpAJtRJAp1//yI
IRdJvt9yAVoWPf5DFmcZAyIEWY+7Cltk0lu7kUkNEJ/RA3XQIhENljW8O+U94wJjmuy8M6Vljh3E
xgGV+Lj146h+bOLr3IiAqz6Sg5o4K8mA2igf9PDBZlsL8rS+FnX6E1d60fyasYbOlI1pk7GJkOSp
XCNCph35V+MNwhWlGWeABAsE9xVaIW1i/W2XMmvHE7udGQA5Mj/u6oOq2odav7UrZHfPkpSNnrJ/
3mz9mhkqNUMIuZ+VWCvCtCYCzFzxii6t/vo2r2e93Dg9clQ2VfM2osZZirJtWt0RpDee70qpy2uh
dQlVJTut+JhUCTWwtdFVzpnLQb/DJzVfOpVaOwkCEW6pEZ+afSXyZyQepKiXDdumdEx1OB4faERX
8zEA3GCOTHxjCrAHBfAoGG23EZBFWnUI7teJssl4bDG6e/TY24RusRdSg9voFT7X6XAwoQIqTHqk
BR70RdySioHFFRj8t2z6iPIPLcdg0W+4VRTVrDTN4z+8pnUFSLZTHasWlQs7zjz8i0iLFuFtxc3Y
gAisREPcaZkl7KG2U8e/QxW3W4T83XiPxqmzlR9/A3PB2ZV3iCw2adC2fCtbIzGS5UNhTMoW7xfT
Ui25mh+Q3LVJoW9/7zMmko522lemoO29355bJQoLUeFrLx8Amu3ZZ22WLxs2hKk+uPVPKQj1YB8c
lmDIojxu0QBxiYOxx8vTa8DiVaIKFo+nT5t8XaMCNsGpwA7oHVJo9aEVxNLoG6wC7fa5MjWwP24h
BGiNr5OZX9v6J1G+WU1En+C3GohEAe8YMbAcZShb39XNYZyVP1YDwcV7ftrA6avaqkSHDYES7CPk
zydd/uYDVlgxCjYpnwFdFM0nl5BICs7XZ8g/Ys/cB+lKMGxkS7WeHxWhEzsUIRoxyFU3jVh9biHC
nJHq+J0Qw48z72kGqmEhhZiUfikCkMngt+ENlmE7GpZB3D6s4Ax60bJybE5XN3vMTj3s5g5IZJtc
EYr0h1B3s3q3DdY88gxq3j74Egv5k+TxHZLvarG+3fjghQdTOeypVZoVpniOF78Glvs8+7ehDkMM
IAQlvoqaYLwhALwr6j5Hdp8sIT1lzH7tlDCyJ7qNSpenL5wFPOrOuwetf3c8HaJzugmWw4oMXdE6
b8IN2W912xq0HUHrf2H9mtbUtWIY/0r/m7TocWrsh2jXw2foY3F1sBLIlXmxJ4vhID6F9oHl8JyI
3rY8BOomq446Rc9Nj3ndlW397Wi5sr4qrhSwbK/ClJl5R9HkWlrOuW1/js/hPenHw+ql6QU5dfbj
H+PSn7xEVsTT4G2Dhew8Fjq2iYLwQD1PftC22bK8mOAaKtmCI7VIcduQ/Y9LXYON8jDkoUhWVvPb
kfaO/LPGz+zWgM4Em5ykaEjwZvXzPFDOCs1L5FosTeKflI2L/A+b7gSJ8JKlHxvK9n1OY3PfjhHK
cympuoBujcGkJnzvRuoGxjPju9hG0Z1MrNFwOhz+hzSm9Uq06GTf5QjBR8ORnVGHxSj/qDJKmvwF
mCSaL1JxmIrBkizJsTljtYgFvlYyrNOKVQDsqZaO7P85OSLZ8itYBvB0PdTYdYBz9Qif0pdWGN0x
neObqFFVJUpcmuCjONB7cikkYYEMrdaOQiduCAOhZ4H/6Ued0zQzr9l/9DJSNlwLVYuViZrUT7nH
9tQZKmy8UTzOG8GIY+Q8VnZV/6kcWLs2BYdx9Kn7JeGJsTbcbebB6qQ0u4n1ccRF1F2cDBtW0Tw0
ovTVF8P0uldYY87xZodO9DVE92KsLoQVJSTXw7t8mMjxXSfVLf4qlq8JlVX7CE6i23oa4wIDmp8E
YCG3cVWo0gepYwjaNAsBePn8iKYQ2mkgHXe6R0nVkLgnp9dOQriJXDymkCAhWsky4b0Iqj6Y8xt6
RBK+ubBh779AYvua5uLtXzjpIMp8sjYX8SCIHqrjJ4zZwExKc5FSpFEpmue2c+GZS9BZWnzP/qVN
R5aS0bkp8j8W+S1Tq7ZtZ1I1jAaTpYuaLABCMtQLArvZ26bUDbP0QOj+1OCBKK38g2Mdz03ySXng
yeE7d0oDDohz4BDpdRVRm140phsNRCbo7YJEltyeVA1NrHAOuYZR+ygPwmhn55jRQ4yh69Nugw6O
adM8Vs+19E6YSrx418azCQ69LKSAPz7PMq0k8k8H+mJpvToNvwzLyFrgi+PpFPlAt7epmWkft5g0
XKqbSzd86oPB6xUkHH1csFfEYrCrudYtI5hPWWc28v/qm0ATPG4jiGHPyQJFGx5GhbOLfr7tec1d
p71qeJwM3EBGGRvZEE979Si6Sw8ZnZ2EEKEUXAdSUjdslol6/Ho2m6x7Jx+hem3HlMGTIcMcJ2bg
xjpvFlrt1cGcCAVP3QLZfpG8T3CfHd/7ypOeCQ5aBrIvwXG8ZVaEz6ueD/Co1oig/ozgo470pSG9
MpPtgwPq6ZPpxR0N22wT7m+6om6OhbLkbqoYrdX8SR5/CV3e4bzepl2dcEGMqcraoBbnhJMQxWG7
jgBRIb5JwDXO4xhLK+EBNd9ZM3TYXVrUe5dSOHl5IYzEd7djMOtGT7BQ9TBO20zog/kFr9INMXOK
XM4CfJt0eJfcnK05j+7W1XlmGJMztNApvzBXDKcjNs/OjLvVkp+x6E5DhUvlLGNQC6CKJYkEErza
UkRWfqU3ijHpop9STplCrZiTriU9xNzMlyPWi14lFqIPvrDJKIhSE1f5Td6R19OyywSyDrX7LB9Z
sxDurJX8lHwUscts+NBomXlPU8WOAQNoyOLF9mqgE6Nxcduudxtng5V7KVlsaU5jMr4+iEDX0Hqc
qUxAz3JWfr5JVFc2WiZBroMk1VCqMVVQxspiy3kHjDv9pcInSYjwirPZhho1gZjEq6iZB7ZWqPEj
RetzULyxkjf6lArhp12VIz+N6YcTzBhDmtcKa8CQ5j1XWQUMzYEsfWxU2DOUhIo+iWjCirgG9RQv
ZMA2FQT0CHWEVm0I3t6UI1/HA69/hZpqRsYCYFTI2XpjfpiZRrW5rtpc+S05+Wx/kuOVUwCtU90o
Xs19yzImJQjlU7966At+KLiO73N6I47oIreAinPmB+3X0CbTTbp7JQIMTTLlpCUrMXZJcl7ZZ1Co
WMNWPQqyN9UkMPlHEGLwJFI7TFcAZ1X+U2pSWlSH+TdpWYq+a1Wt+szY5Mt2xfZ9BMcvUeM9Q/RW
Ju2N7YgkDw9smBpi8dGbGip0fO6LQIjzcBlIVQdxkpY/BMDUtZV/tOPTVGZGHsphuP68/1UfdfYh
o+urUq1A3gb0MC+BIxIVBvh/KqXfYngzsDm7VQlGPOLhR9gjDQQS0El21JIk3keiXmZNF05Is9JT
P45UVwEB5XFxtz0Om2mbpbBFwFcx2qc5SeuU4oeP8pktAdjC6BF1/evOF93ebbNCBE58EH3NoBMC
uxMk5+kwSTzmA593dGynTkOvCS3iL2qoAftYijASy0nfWzZAZzgLJ1eBpNdjxASDkXcnDrq3JXZS
7dK3w7v1BLYc7hSe8C7y1InelrdOuiZNwfQLCmUbD7xInmRwWAthjHmbnudMEmK+aBnJK2MlUBDt
5ifxnfFaRXPJBowBF/H4WzWJs+neGGaTWe1R8dkKC1xRkICso5FOe/ChrvgChzC6qWAfDW7k9pug
aejBpFmjGybQxCb89rZ8zZJE68/A1hgZKT645pBVFxmxFp5nJtAZ27OtBrQGJ+8i+okUkti0mgYd
vlKWbZMNn1vZEe94LTl6ZG8saOhDxaGhd/m/ZE+4do9rF6B2gej1f8xRmrQvP6HBsaDqwTRMsY70
Mbf0fhgDErm+TVWSiPu+bXMhxTk1LTIq6OFrQe3XZQRByf3sODeZdjV1skEyIZOmzFRj5axF6Ca8
sFVWk5qRiHON1PjaNmb/uOM8K3+DlNat9PFl9LhDni/Sy1hptvrVl+16TEpirgTJMjVAk4EA/xz2
VGVwm2Nxdya5GOoO2yAyr74/H+wuqObqVwohOPKCF3qgyvfAhR/vsbHjPiKz8u4WikSjP44CEjeV
OMASW10Kd9kicOcMR+j6n2eysKaHSASdOcBVD3MKEuTg5HNCXfAcTww9TSROELLy+N56uvz3xZtT
AhERxQKYQA9NFz1NGS5kKrFY4b+YVS3sG9hMXjIS0RlIR2WTDbhkjy0qHlxhb0qAd1+oBFXsC/W0
Zh4McWgs8vOSyHNa71WJa/puVg/fCMlHfOKPRtaec+XKDj8BoT9FSJZ3CJ+3kzjhJyNaTgW2mAAk
W2wonuKmZXkgmsb+I3jb0A30KxJ764KOos/UtoWhxNrjWTPGgrGuiZz8DyFIOzLvg8o1QmUk4d+f
UXEe9E/GrjjGj7kmcqs4RdAJgQxYVdjkk6o5AQE3aC3yiJKDYgIXPG1Oxw8jph0FLakCmg1Oga3w
ul3JxW2sV/OhPmbgYClSsXePTWgZne+VSI8mk4b9YkDF2SvKlOjtwooTT+XTHO72UzBJHzrFdeLp
0wfD6uEWCrT/vESZGUZo3dT+YgSxyUyDuMh1gS6ODsa35HinqkkZPldmMbQCGfQEYK8UbcSd4aBY
zbtaLaydcF/5UoK0E/NL4gDsO8YILiBpqvhNsDUSxJx4jqBABhGDw6kvEadFaqBbxXK9uR5/INQT
nymPUYNbIyGmLoitXZ/xwZdaaFKIEMAAg/CR8go4EiOxbUzHTVBeyQ1b6KmnCfVwa4yqtFuH7h0+
5AdzK1FCqnKVDCXe0+deV+nLxSoH0hAWHnzIpejE+taCs7z7GYiJhcDNiC6KaLysgXH+dmY+QnZh
IPtusnA3oh0blXIvnZ/bd3G/p3ERbO1N3YSeBCMsRlBrZgIGEdtj0crdv7/eJn1Z7huGDZext4Hn
bhiBgjo72SJV1crW33W5UzPUWCu0prk7RF4iUM+MdWUdVlDE3qpftQTr10+8JLWpkyCFgxpvyUmL
ms4CLU8Zm131RxLiCaFhcyPPF4K8bCUmTV0KemF+VaY4dGxaEIOtGHcX7gV1ZeaNyOilQ5UoseJv
ktN5NsiUYL/5KdsODAxeNypX4z/CW6vzzjJjaP77sk72TjNJGeZs/+r7GuQbaudtI6HqCbJezebB
lNYYyHlOtmY6RJAC1p/hMTKksBpTEefmFZormgE4tIAFrJuulaXsQf8PTZ96KeLZHW+Pjhn9/Oi1
2TmlcHVVGAQJLncDy+3jqvGhuncimnWUg5NuzO1vkrFUhaz0aEokPEDBicQmrne1Yau3ED+FOGWs
gj3+HZTjtsCpWLNe3oXwW/Wu+Eaf5Fz5aY6PNZgKhDUZGXJRHaIST4/jcYPawBzPXbJhzZKtjh0q
at1y9blLeBcx8aRVcVXBsD7+qJiHErhXH3HwhuG3KnyP7ZS29MAmaOGaEVw405Ojjgergkt0Uuo7
TnJGOpvpa7Qy0yscZiv4YeCY3OVla7mTHgHWk8wnyIfNn9j1KxoKy+xv4kapAzYja+4M8h3RXMps
ljlWPQa5q5eec5gJQMETaqVYOQkducocqpqIGRbZ86F+DZDb0vZDw0RVhOS+XXuIN4pkPoDAakYL
NkHTZha1aUaUd4RS5CelWUWRqh7NMijO2ciSBUAKOGgKVqeoVfByJDmxRpoleT0irf+G0ACEUsej
Fo7K+OHroNmoEopK1iXS71+3xrJK55AOxbRlQ4/c74vq7fc4rqRq5gkTt2wuoj5TdpOa71tRXeIM
g8XnIiobMmy3XUh6IW0VACiT9oJjqDBu1ri81sKa+jUwML+bYsN4va0UCd+scMtEW5YudY9r6CGq
PHnArRPx2j/5uq9U/uY980jt9wNugZpnS6/OPkHseH5EEG1xH/49pn7uax/HiLximo7RKGSgWkTY
GbuN/H5DqTatjooggoUWdGwJDS8BBmVGUUqmGn4fhE2eVocovfEIAPfcTc/iyXmX/XbwbJlesSFZ
T35ag5N7NwoSD+o1Ea1IDZxRHNCkuderSd8Sxdr0nRUsGWNkpJjjbZj5C+qfCkeqrf1KqKzUYlq9
lGXcRN0F8vtHAc2QOphNvy3TP57ExgFkuI9Y4caUQHsErjSBsnwvXH/p/5gSxhLTJ+Sx3Cy2+v+r
0gI7IqXbmYEQ2lBI/WCG238NE4R9ZYeSnPzsaZK2hS6jktfOHgwcD6Ka3mg5LoalXxKH2JfdcxeX
Ti6WMyoqhXL52q31fjJC5JqAi7dNLT+PEALPelNHZHHGFY+FcE6rbmajDh+uev82kGKRuxRWe1f/
twXbjZNSMOXhWyRr+waikPprGFlFaqBLUI7qpJjwwTgRSSAjcNAkyWoceQEzjs1hfZ7ziCvZoDtI
5+lMdoBPMCg+71qYLOp8LiqBRWXo43pnYBAZiZU5Sq0O3f7cV1g4ipMMTdyS4DP07odTVATv89Dn
ok5S+DoH55VuNrB9lnOwY8bzsPt6mFz8MQQnwyGL050C5sSRQEtIe6k+QV953JCYnL/FiNwLaDJ8
ynROqys51VwoOnooTcYl0yjBhD3fvSaEXeY7RMmbZOp7Ig//Gn4KUoF5+LcFigQ1Xo1yo56MfH3H
UR0W1MU9SB8JnDHnolyTMTIC6QeyZNgbsYGpUpR7jbIqI4+Cr1Ux/Qb7xVtJcDehCMB+r6DgAsjM
nORgl49E9tOl5e//htsXWhbMtdY+ewdTtnUICQUgH63wnvLQOP+gG9gqqo3R7sfc1p9GUISc39Tx
ouGJ9J392rsxa8kwxfDfDR2YTWp1lTe6F0bSuGyE0uLv/TCO3TqrG8aL5/LAR07RH3LY+ObmYpYI
DcAfitbt8VgdX/4p696V31H7+A7IcKRpk6UfDAeAzQbMo6FKAKLPp0JC4s6ZmSyCQvKo8juFe3yT
tUXD/YqfMAjUYwpZb/+UFLaPXoewVUn7hooFANALbwcVWFgegLkpNHz7iuW8oc1jbXyL9dMrrqqv
Qqdob2lmZ2YhceFWorR9mWdtSNCsTFn7Dty3CiPWueubJD55WQFtsS50gqQVDfVjKYpUwMYYFzSe
lbtyBtUUwPrUoNq36m8LhxnRyylCAC7vkQTFamglIkebVpkVDALfAkFkRt9da86G94CBDNBTWjvQ
KLsXjsWkWs1oiAhiuSoGul/PWGV3jpR7KV2B5CD9qbnaqUTtTaoJIFnQV+yEYZDPjvugckWxJfPh
fgsIzlgwvqT54FHbsx77ilNjCR2LkqtWivl21L5dtG0NYIbnrRrNjyN6I/ks4+0nZfqPG1jpkhGy
P2HLmB4oNX3LkSN+r1poZUM5IpSqw+Gr1Cp1cYzGcpi9x6gaPTndjBJcUGxh6ZiLuX7LiDvTIpDA
iUuhHBUTEo1CF7KblYdt7iJV1AmmugeTx0/vMdPHSNwozq+HNppYwMyfDUcgxIRahhNKMhRoIsvQ
PYgLyAchLVtQuA1ERe75p3kuzXj1chqpvGDjIcoprldH44BBo0EReKreHfeBqZVH/yueeGyflOkb
3ht0Xzx7Ip9XmON+iQMwOx9RQffiRBqyi6PVcPdM6WuG2T21uy86x3THwf4Bv/oGrfQeIFzYV4nh
2dbbxFoYmpuK1JV3FFt6zPLU1B+IsWNrGhT7C9dus/9TTn8A3ccMsntSFTg36KKKvAK4gsQge0ak
Dq/5Ki/Yr7OSzd4x/zLg7XXs3GJN/nIhX8Kuom1nPyL8dtmwQ8lQ8lwVYZGsPvUOVqx3CpsRu5In
qyQB95fvetAGlmxUzVH162+KjlVHU9OTOg2rJvg/ggBTwxPczLkEONvUsPNTwzCNzYx9d0X3idow
t7w5F7OIi906/fBzOaUNOmUXr5xRA9IRPXVdxSsmArX0NF++BDCbLt9thNZ6rJm4VI2vHki7K8Mq
T2Vi/LzC9UO5VcbOcT4J3+g+7EaeSuw8SZ1S0z2aDDSp/YbujobZL5YwaHKpQPJLm/h5ZIP28756
4xa4TlioNPKmrD0vf+uQaDNONTMQcmS7HWrPZGNDvaCH//gCe3L8Zygf+Jxkg09F8Eutpa7tgmw2
7fCPl6UYHBv4kcU6NLDn8qRZnrXib+VJaUBKrJ2xJPdJm8WhnOnqJ8FYXzFraDnq2jbKCcgQU0bY
rmg52Q89n+qm43HZz82O9idlyk5NOo934+tIMUQ/QfwDOukLa3q0+CDxPfQ4+bWG1HhNxNLGVVTw
EfjX/stFSADYARTyN+8q8KxNxf/MSj9jo6dCrcBIXn+kc6sz4VARNprEMczYaWp6i3vEl68xY2uU
VCzPkg6safW7Vh/WTXbKMi+gDQrQ/NODVzC5jetSZLaftE21897K23ftcKf9/7P+QIErBj72bsiE
1vTM182Fwpf13ym56tGq+cOgWJ1rX5J++bXFAiUytbocialFM1rJcVWmUFqXTqH03x3Q0vB0b/4o
XoIhQDeLmD0QBv4NmJZKEpLgQoQaseMeZogVml10d7mEx4SVTsPfYWTBmw4ndNdDyzpyDJicYiu5
RZA6HhcQ5u0Q2djGtS9J1Gw+Xo9tk/iZ0LpR8vO7hGRkbRONVdsx9bkStU7eWph1qakxvSRS2TVw
N8NZ7xHzSjyRFN9HFU4qV7n12m0mR6JblK/DX4uI0WIw2V/8qRDt4zt6PsQjchsMFuE1AymWXfbI
YzL7xmrfD6nQJLJrHSnPL/Hq3Ufias47bDUnUPMZ2VdoVmbdge5sK/5CyoVq+q7RQZCmDobBKlap
em4fw0xoHhgXFzktAR67DGCyrgnxE6igoQloLEONsJ96/vLckqrHr0dYDi3ZZsklIEqMym6xViKU
4HiVCiTSafzsqlXn1HZWmMAmRt1K3jj0NKIv6WvdhMgSd5x1tg+cliavQeXP0r8U6XfJLvPDFVRb
oRsfe2/7dhuyNnqeXivjsCT/Fy5D4n038EslK6VQQbrjPaG07kcHy8TWKjQS731GSu7AZAwTzTLJ
m3vdJBGchmqBgaIBD2V4zlFG86FTX1rdBZ/2EkVw/8qE0b/2Q7S/ynAUtuh6O4ZovtfI8+FtXtVK
5pxFtA9LvWYZhNAKY7z7IV6nUHtKJrCMG2f1QAoBDfSfnT5UuMeALMOfJvnBXGs8l7Q/yCqPGOuf
CWZAFjSZo/7WGO9V73NQMrOu8Qc/IkW0x4qqQro4OkSru+mZAzzzBu99jQbdH+WQwYLqirKkPNQc
tdhYRuvYBPODGRJN1ByicJhdXJi10qZ/HUGmu3Ilo1IjGuovtTLdUZknADx8xeylvJRlVGQosixf
1p2xPqm311I7sRusdV/I5yVNbkcdeHxn23TMkV3MRc0XIr+AbE791Po1TWSMNSPdSjc8d3yx9gVv
hjx2BAUXjChA7izvZOlddj+eeuvXeE6PmfMOpQxR3a0fyKbS6AP0sTKmCv34FWUklsJEF/y88TKD
B3k1kFLUu6ov16z3rES+EFpUtMt8zMUY43JYZ5rxCbYeyGoMJB0eZWTXCEk33Hru8quY1k1CGNAQ
zalaB8Cj6yZlDnEPjaZqPEoD+ew6rhRx/KKakFCAeoCSc23wdplD3h6NCNNh+hp8+Rb56isSR4Kw
waR/B2nC/48z9FjlQaFXY1fPxvwkqHHZfqhpQGWetptIqNIf39AwuEKVqu3hmLRoHe5sBFgTrd2U
lNpyacjetDMIb+/kxJ25HYZmSLR4guBcEfJybfOdb239ihkCsSj6ypbPVpVPTaOHahQ9MbvfGYSi
oCD5+keXEJZtdOiwOkcmLBddMm4o2yrpmkV1C8XBf1KjrI38+IUapyT9Hbs0TSDMMESKbsD7dzkd
rS/edEZhode4zm/SMqbY6XtoXpiSfUWa0lBbaHHffo0na1Yb4ijqfgvIbjVL9pn5INRjLdCNUJLP
h+YAcWSkU1ADtm8cV49TYRgLbytcUtU9LLqKZcTmKRHYkmt7fDmtvHKcXXYk6oOreBpUxNz1YCyA
DVlyxgYn76J/7X7oumIUoQeArTs6gvAXlTQP3xFvhJYb/YeM6vq9OGV49fZMzbbusYNjaUGgL+qv
zgK8zb6K7pA0RAQP223ojqN6Y6WdKvuT2qztkC94tbV/m/yRQM0wl2ZuviHqnm2+rQDL0xOzxSrV
nVvaak5HRaNZczqzy1KwoPBic01qsPWhyzvIwT1TCeG/8x99+CxZ8nflreSZtXAhMFTn2KuiAsjM
U+qK5EIZT1qXiuwWiAgaelOdLwu9jd28B2r1Z1dxmjyhN72nCWTZDuYCXB5jAJjTtCTivQp3NoZ5
6/DJQB/LkjdWunC7uRxUsjnW6QLxhIEQ4LlI6bq9LuEKeEqwWmRxIfsme3cMLmqqLPvwjv1T9YBq
veRndCMmVd+rgvNvXzcj7GMBWz0OeU3eM+NyP0hIYPCTXwOT0MzysgoEbn9Qx5KWvvl+zX7H7rGx
FVmy+1qgDdJQvCk1lYuDwU9R1abaYRNdXN8sJgNzhonpoRi4KE60LzGKjiXOVF4+dLnWbOiyaD9Z
KkHyH0B2CWELZ6EprGBoYmrVVDUFy/UzsZCFRthzxM1hTR8a4nUYiYmnKUfERGOopXERRhIS4oVr
r3yZtQ8Om5KZAwtXXCsZpJ6/sjiojSFsAFvRmURSuDDQ7AuIWXCRDmstxoY1FzEar7CuEB3Pt7UJ
BBfiV+EU+bw8bcOAoydX3d35HGZ80fyJmAedJ9z2AS1YsK+5DFS29Xyq8fYvxeznjWvWzgslGnkp
IypsapfT575hdmr+4mrQWh0nQ/ZlfMctpYk9n84MzLXz4fsBqzq4wbJqL8NwI5tB2GdW3IlLDDoS
mR8cn/RPWw47p7lqP3+/F2eNqGyAZdt018vS9uLcib80/YN/u5tVfdgU73L7867O29JXmei6hg84
G0x5MVK+SEBF9bZ5p0RDWlXEbYMhKcNexGwU0H03x5UdX39YVDLaNKiQczyKfpeGqe7vvpCy5u9A
mEy2Zne6UIv6QBZhR/A3j8DtnE+ZfctpyB/B9A40yzmGjQUyrOWwyO0twozwoqEO6dMaWOQwDiL9
dAZHuXbhXHnBpWt/b7EOSeegMkUgKzWZjX/hbo+W85dEwMV0Gm8YSMXlKIhcgfBJaNxrK4ezEBC5
HMYXl4sitBYn6ua9KnTPXKZQwn2Jcj+NfKLsnGqaxQgMcTr/FwOFgh9EtZWsAsEA+RhfHRZJQBZT
l9CfeVad0rV54gDMAVtmWaPMMEjQAqdn5oSjm6U2PTwaItkOvwZxLDEMy9gblgd3Fq50otIw3ypE
LIfH3S1PT17qpOx6yyi6Ogu4SkePHOuTsXkbTz41IWBTsXJVQ0gmKqbI6zOYinfc+WgWmE1f9C4j
hLKoG6IGO0TH/9VPNGREa2o1vB4mRiccuTkeVh+pyLFOKSMDGQWkiU+uZXg7/oLeW7JfjB8IakHz
/ZoucF9ckICjvCT5qhj2XPbD3H1X8YA32x62qD1QwdTr90vAHQGzX/Ei4M0tGu8eVGCuqT9No6s5
NFAD5S+YHhI+/2J7d6/l74c2VUTeQYfmpapnoYkN2ef6NxlNQBVeZmh0I+dkjIwJOMVkyM6okFF2
2EtDQ8FiP5IvBFwmxL3YvSXk0nsoNjZG7E9anou7OxRcFqLrpgPy+WO6JQMQJEqKE4w10le6OjHE
XHOZ5rs+XeWk4nhxWK2RoiCBSOKYm4OvFHb8nAPF1VPiWA/abC6zY2xjxhEIOGHEfgB580IYNHfL
UxvL8UOuFeaTXav1Y2HrPriTpu59s6WZKvjR5io1fyGR+p4hpEVdnSivMyYFY9apZqHr7gJZssUd
NEX7C8/G25nlJifTKEVQPHMACXWPEzNqC5UX5gJ6303NlAJOBhGTguw4CD/xTloDx7ADI37rmJZo
qoGoYHkRSnK7EZ6ZklX2i1h3ZcqG3m+IbEqUcptTUZysn1lvTPgb8Y0OK9eKgTMOcZHIqPuLDmky
fh+Nx62zosQKkhGGvxrhRyvSG28dI5G2PQDGMBgRLRRg41KiMTvJswp3mT87JWychT2JexyLjj+s
F6uL8XXhi7Rc/5A6t6qoFAh+4pnRmPkrIT+oGk53PCZjrQQ1bvCidvI/B/ysCgobucO7Hbv72ZX4
8Lks8eMCfe9+5jijEHdFg6goTBClhuuHxtrENY/cU9M6vATrHUQu7VxN81TpLrYum/bEKekV9i/T
SoqrTW4Zm5AbITxDG4vgmejKcvpNLLQ4IHISQuyE3rvfII494jfP3LrDVemhT+XMCcCgnQ/tXzAY
wJld9F/vHd2tq746donTaovkJBpTemSQ1s4JgiU5STPwBcTqS1Yx77j5vRKTnaRx/TotNvv9c/z/
fRlBhw8I1zHuIJA6b289wMfjUywMESQ+K+ljIkjmJy7pnp5OlEe/aLec3eDTHUuakdsFht3ZiLKk
16r4ZDNwA44vgadFYqt5njz04odU1sKZfCYuYEs4RW+6tsno8C9pcNvBwyLiggsRToc2BHUH1K5T
MxIN8EKQlWYUSCsVR3VdI1TCh9NLMTx+lG0/MIsbU8bRJ2DwvGwW+0xZ7RGb4Fq3Zg044XVGKaih
MhsLq2YjHMTKsH6eV362l57KuRi4LKGQjSlkSUyMeyxu1wv6/k9cmGFtwJ1ktrCYzdUwWLqhc6O3
yQodeFrakeN9J3CrHvC/ewAAeWzRyNtIvsui3008y/o0iudd6vPsn5grYOo1X8YXoffUH4I40ob3
l9dSE40ISZdoqclGCR72ZijvzxYmMbZ3n9cqWonvxzc8l7XSNOJYKjNymxK9N6Lvjye/z2SRNLXf
NZy9rd7TPjg914av53RelqIXS2812peGsIf/IBOlAJlaJZ/SbsRZr0hHeuM5bqqWd+uZnuwBkjMd
Ls7Di75F1pUJd0zaefgwHouCECQjpj3GzpYevpbHh4YEyHK66WK1d89pR1eqYRheYxTisHFWEtY3
IsvlR9LZejIIMlNFNQ9wuNidiyST/2RCeSctYAjnCl7EY2ayuIMqk8XvB0cJR9BRERO8lwKlm0Z6
GMYn1e5QeKZpg1xnrPLLIVY9bsQvgOd2n1U4ip9xndtoeyiTMNAOL7MjegKv/EnlndpEYnPudWmb
c8IKd3G28qwAJ6Z3TrecAhUGy8V+xHJ/OfskjKoUcu4O/S/+PnI77+Bt5APYpFNxqwnVHSHqLSv9
XmgCasHFunv2dGt4+rXX2Gb4osbR4B2P4u7Z+Zp10Fm8ALwsLu8cKdfm1lPwlloE8bOlxqEcJWQh
zKVi0lh/HmopEhUiUkzeQ1evEVjEMI4n2+B7Ol9E00UZPtHYhc8vogSmJL1dML7k1IT0CtfTfEQu
xDaLux3oSOEeL7LHqeL5YBZ4pVcGUGcsww+2hkIkOnzPjfE+HA5VLDf5vZPNJ+2oukld+1Lj6MjU
ZjZ/n9mdWtd/Sbv4evfGN2+J2jFIFnuVcboEI2fNsJs692O78wxfLiD6+jk+kOZOeTg9ZFguCEch
OKNwmE0Fb5Szvz8KkPYL1jOt2b5/tdrOqw8qCntbr/+nomC/43t8Ynz0+7sMEIrM9Wr5ryp+WOPm
6K+oI1wBmmS3T+bjx0Ybn29k6nglYkahasY+pcN1z0prk/0lJR/WgqfHOGCSnXorxRZhs98VsncD
S29ECpPHEP12twXD8w3CGa72++TGQanQ4npqqgx51cPusmbCb9tpnGUS5bkZOsEbxAVaIuoeviDh
qoHd0lnmTKFdIbVD/AJ/t8rXskGGqf47S2kIAUggaO9MwtqkeSkQMIdANuwTDxM47Rio0V9dVsgo
hbq5QpWYhuLq7jOFtcEhudJYeJUzVvouxAsBnJ5G4FZ1kKHcuIQUoG+h+CiD7Q3aDdirDw4BusiF
rAujV3Ox0N0cZQgDbSOrOcAUVQYz5l+PiHkaOlVL17IIxsfr15uMCv1CxtsIXafJ3Z90FYDTava2
uzU08ZGxmaNNdwlD4UcfinrytsrsxH58Bdza7t7PCF09iFAcu3MfnifHRfnYy0mfOS9KSarwx4UA
kiYMJ3AvNGzO4cRnyZiH6/H9Hd4oQLu1s9N656dy+UW8Yu1jT+jiwWxIujcTwpTnlWDBnRBgV6Lt
Se5AWoF8Q4HRqAkUHPqov95XX+BZZjYN8WfNbKKyT9dEB9LpNESSisrbTNpgjxiFCh78whftAzxZ
TKn0XFijRfUQRFHbDcUSnDPyx0GvMrQzZDbQmuGMuI2gvmctJ5l7WoEWyEdfKkfagnGdIGrbDzKX
idHl7lPpZLbWuNsSzxtN19TNh8ia4ufnC0sAIMnqvvDH7kSllGpxm3y7y0vUofi5u08IqS+Lp2UN
dTZf7cDKn6KDMPBRteOwkTgMpc4uRhSgXUPYDvB9FVXVyt3iR+Gd1TGlHFvULdlrrE7l1pMcHPhl
Ht8t8Q2mPFqXNnayZpFoDKCREnhgasDdTmDuhKAoZCkCNOcu6CD4WJW72FzWwcT7GiETQ4KBJR6d
TJr2u/BEBOF+lwE5rck1KpwYqW/aCNPFw3Rmi0m63AxQSTu/FC72eHLOQUJEKRUFCWYYkgX3c2eN
/T7HFIFlATtxaVPdSNVbq/QM2sQ0YyTjuOP0FQWGYBIjJfuRMSikGPr6+SP/0VyYDTpJslA7Cox2
QuKHUISfo9u/dQqJtFIYO9cHtwEPXa46SPJdZ8f7sd55HwjIOT3DFiR3zHPe9paA70PxO2KYrm6V
Hj6PqqHjxpIOg47ejoaMrUlfpZ6nautOwYgkZ7GlsVcNnHpzCiE+1zjpT/sXlcrFR/Uh/sdse+Km
g3BKD7HTOtg93lnZUYmVFXDkyfyKeo5xhM1J6EwoB052v9+a8aQUMS89hF66Jlx+A2xPuq0t6ovy
XVzAomXW667VPO7HiYFu1on6r+zh3qsgyC9/kHJmJ46crdk42gWfenxLn1hFm+Ef7xFY0waS1K+b
0G74wfFG9JB3Q2b2LYyGhkGsxMz3OUomzLNuezuu8Guz7JBfHN2jap1NfLQxcWkKlq3EXdWgV0Fk
3z6TnMmNQfgbT7NhdetP9cBD49s6ef+0t63oiZOwWHSQoyorNDKUgE5+TXumBkCPLLKzAQB87II8
HkSnN2J5qXYGpa3SBDenMKB7ZtmGlHEOcU01w1Z3mH3U8ZXe6RBm/HpVzQJLDFi9KiPf6CEfV7Dp
hDfaoZ1+BGqTna/rbzeoLJesKapYTNVe1eKbX7eNADUklmp8d7TGWST2JJo0PSn9wRqFRm7EdFU/
VsY/Ga8LP/SCt6sM3uVRzyXKKTJ+QqP8b9fHeUrU+iLslxM75MqRFpca0VVWd7or4OIuf4mwicmv
wB6h4FcDgtmx5U7GNnvfh/KjhELV7QipHumOJWG95WSxrcz263xDp3b2NvfCcFkEizjI5gNlnTwL
oQs/jNMywWFAXkMKx8MRoKHk+N2Pawom+hdRej3tpC7LEE9OwHxraBgLLAvRuBV79iyNjq/oAUud
j1+VQrF8X6RSOFpB3YMdoBtr6a+dv5wYfpxLxFI6gPe2Vo9QboDgZY2k8J+1gsIEMeuOsqy+FNu2
DEjGc/MzjlRxHGY5j2qT8ctxL50KHQ8PJcSJnxrd2y1h5YEb5l2ylxVD87/ojPxDA7TuBrpuR0sf
kQNa08UOiEgZkBg5bRJrA8UP/njmjZPLE4b2aVLQaJukoC1ANgOqlQBuYADFuFIucdudtdjlc6r3
iBnKCRrPQxD1/digQ0GT1rUWywCbQgU3HDKbTpNNl4I1yu4/k03Lojo4F9Psflm3GMhPX335kyNu
DR1OGvrqwntOwDwA1yrAtm9+5vc9InGJF96D/Lm4r/CItX2Ht5TpPebjrNpaOMxdbrxlm8AanAsm
eYJOXh0AitXGOr0CmsdsYyJTSAm99KZkpo8XKFR6jd1+UV2oQnniZ5BLNEDSDyD7tN57Sw5Na4tj
CHNoSQwpr91byJ3PYkmuTv6gIho0adowhPU/xjEoPNXC0mWLn3M70WyghKM0pBeyNrOudnIyhLT0
y3QxK8FQHJXER221anq4U2zVRHy+OmhBMu88Nfi0dNfBvQ24QFlMx4ORSDJ5zUtraLwSF0ZxD9qP
w/ZwcL3cfXXXNSIKW0kiZbPFhOKrIWcnATv6ThSlE62YuHuMVXB7ehTl8KnGjD3ELQsZ7IFDA6u+
9b7TLTCuQhRLryr9OiUXNDAvI0skknPXTxLmyh7WdX1Ep3EOdnKoF0J8yKrDHabIB/jDNUoZF5Fg
JJ7lIk2Hb5IPL8jo1y/OR2XB66JWMAa5xdjkGNAaV2IkQVv88Sn64sB+BvCscZzQeHMhquHtogeX
ZjQGN6reK4JFnQoVKjwyHxUOq/10ccM23eLEgKGNo57EyGYqFl2Svqk9N1J5AlgXHwu+OjzFIRS+
NcfuI3RZZudxdMRE8y8KnNMDg+Aq27qH0d+0SbVNPRfLWM4B7qcjvPgU67snmp8FpUTVVshh7kEb
+mGMlKpHacaleNaiQWIJZ1drmpHevj9QJwLfdxrK2BHqXiLCe6zWXn+OYNryrH6z/JFmmMGUO6xl
G46qIepy+LJk2df7Ft1nTPeZ5to7Tuh/QBkHshRVIYEwrwTwbgnBPV/+D/1MkAiwVr9PO341fhj5
JVJabkWVVN9bdeA0wtNnYiluX77Nn3RSI6n2+QniuVTkh5twpEx3lAwWWuAsRp0u2j2aGW7kYtph
qVJrlDG5mnNxOVWuNjRzWkdaQSHFcVevhywKMj53jVydzyl16+TbhALPyek33Uu2+BGTqqbz9Bns
Wo9q76BNlcdjv9nRDzZuuc08qhy7/wdpac29cayyke9wOgtJ+/k53LegwRimVol7XC6CVPc6w7PH
XvQe2Z9zQTBIsnlsaiiqYoxfpRfVW2im08RzZdWPorKkfR1kIhQnBoxmd0HyC6o0fXcXW3y750F3
vT2QAg7Nv7/6ztbydSPUYb53opf3FymtoPFBrc1qpL2/d/JFAGNyKGZadoyLBvj14wsPMvfaMAlU
g4oQ/mYCfPjmN5tE1Qy+wqF5aNnDRUqTzhRhbl5uK0nQclKkiqbrFHAuSCjgvN4a96NFbu7Teo99
Tr/vlKNZ/VGyYTqFvjRHD92Wv4MBj/7uOrI8tgzV4qHpuoMUPfILLXSHfE0eDHkeBBfyHO8bYBq1
AxkizIPd9q4bh3CQyHlSV251+0fbshq9HosROz/ueCwGm4GS56GzYZXQDLdcZujZE8mYRIxiPkfp
iJbzdvSMwQONgAPVgsyB3J8sZbRFkQNYTI1UMAXDGBIhr0GgKhLwL3dE4zNKYA3f6Dckn+7yP8o5
qPZTYJW/MFuoNYVT0rb9oX1a3qxLwOvgVWb2JYdwBBdpny7Zlyyilu7ggak0i1i+L8TzQ2zI31YO
CL5f6CFLBOoFmou2AqkACjPSseQY8WCojaE3f4Dnas4dr/7GW+XrojQmO24CE1omtJEru7Q+7KZY
YBYZOFCKwM5AgZR8HwNanBufn9EEesVcHIyXQc9v78eVNnwhLWGcc6h/DGRb4rjrdsqIuXFT4kUq
0e8jLkjoVq/mp1WMbk9sCXrbwp+KU8jlVSiVLcQwcBaKLzbc4Zw+KnV8wGrRe92PxgJ0rhXvDsiS
5AV2kE9crr5AVBPsaFtsTyXEA5fHIy96TPifWtTd0UzHfca5azqkKOdKobOVS1R28LsmbnRau8X9
umMaJA4iB6kpu7L/3fD637cyGe36R5lY9BRvHHobyUOulj9uaOgmFqW0tHtZAONd5kN/kjDxwyEK
esvv6Qn5gUTUZ+M5PUeafI5utpaxfFiqEHfsElCD/le+g0x7+iwr89hXIczK7Pi2u8DDfDmr0k5f
QdTUbLyaWZgM0ah/MsG4CBzyACwiyHBawCvqvqm7pUMFLxV0XCRePY+ymp+6I7vSsC+9AgswLbTA
F+kWZC1DF49KeNm8NntphAGYTfTac0ApSPrsrjPf+Y6vHD0crw81KMKIn854HqZwJWAXNTF+tNDL
GKB09mtRPABfQ66stUCEDSn/wk+0EnLS5ssugIHruO+ijheEwwPaOpkEYO5bXb8MgSjyI4xepM/p
AZ+cQWatVy9CLj0DZ6I8mNt/Rfqch4qKs2hVpprWbBoh22MA2a3gCO7HEWG+aMZpFR8hjgnvplcz
AG0FfKUJ9M34Sktk+P6KU4xhONl11jWrlTvaMRvi9N3Bc338qndQ3e+wed/kfGMjl+kfDvzR7ufT
1xddLeMp+4oo8baR+iIyvs4Hg9uL+8/xJohMmocaMFvJ51xMh8BbSxM0cgpsmJtowF8CzyPXLXFP
rPklkofptksPqKzXywWGHgNUgcZ/GdHn+fuQZzenmNAQCwUsEPUCcgWvP+4yDyz6urdMPmVseb7i
w6mJB8Odzzoo+ppx+yH0+CgKYy7G0M24x0u1NaQY+hqqEmk3Fag4zhWmqoR3EKz0XltZ8gqvj8gb
WR+B/LUZ29KgRBZwfLIml1J7tDkR31Y8jHFYoTGKlh5iSUTkZDnTQmsdom1sJxCufyQYN35u5uqq
/e49eSvlVD405c2N/b+3cgJ7N8QZqj3k0Skip5tsC8jNURkCcK6hNsca3gxkrrH7fZvBlTmpDLho
IBkCvomDykNtHA1/RZ3+acO0xvH81powJLx/0ZfjF42gkplx+K3nvylekywVekcpnVnmq9tTstWB
r+ta16dlDLua+75YzBila6bx608lddhPfqlYBznpY6MjYdfgei58sitMe1U4unF2v5AyzErNSx2E
vhGUgBkD7EbUb/KIi8/hgIRpK0BRo3VgRLkVHfssX8iO6H9ha5TFwcxb34JhF3VZ6TuEggJZovLW
+6NHPh5DjiPeaWInmEp42jB0/tX7rFqplDQuocEM/O5VfckYY4ct0rwBCA1buqqzZvwSCgvG4MF6
GPoDkvVfWI7Lf7NjHMbFX5Pu8ER+wfNzDWP0tT7ZkU2EjdUU9rsjXFygeTwAzy34+VKt7WcIo0oR
pnru0kVZqfi7JcdsNSXFwihyyquU+DdcLtzqbkvC7wBmSCL67A2NA/dS4+2zE55RSe84PpwOfWO0
UyEwoyIG7G8wZ9j9HXeU2UWPhQka7f5Gft+ECtPxQy5DETOuD1j+06qcD99ugKN+qq1urSRKdJ0Y
yjmlG9sGaGlCXS8be06rsdHkEetYqgFlK3kR5eOA7vdqKaeZgl1085dCVhRxQ3AUAfLDLEqPfaQr
R28XhdyZjVMSVzn5Ff032p981NE6HD1r9D650anqEOFxCLoHHgfN2uYGv/bfWyE3JRSbkg92jjjB
1fbPfDCaG4I4t9/twI2/1PR3ZtUJHzHicjNY4hg9rTn9gwoOyBXsUfj4bfXzIV9JiT+kXWFYFfZA
AcXU7wB/e4+gilp3Z7IHquWNU14NEv/3EQuKS/xgXud/oaE0KjfXyjIkr5ZR/4N6Qxb+H6yp11C2
1VtnjgTqF/v/oCHJM9HvNbdJetbMlkk0kFvu6jqjKKZZXfp/xxVX0oyFht9oILLG5olGoH/l7G4T
uYyk/93CtTQbfOVn8YN+sagWcDmuAb2qr5bABNy2UF01uB1GDhBKFALx+n98PHqCT/C6yOnzTgVo
6sH8vXVAn3DzkIL7Pb4Y4Sx4D6T7TMdzru5jq+U5ZBpQt9022bxkmieyuP3oMXU9K3FHgGphrKCY
o48XrfTVp0WTX/UUaRQEITXt+3WcMK6xZdBQfVy/nwkY4OqvEMrLIewCaS6fiNUP89W7/2hgvwrK
vIrTxdyyNSc8gdP+DqizhsuJrxGNCTlQy1GFRJffewkyphpEysNwl/wizIO/8fj1hSjvhmy/4TTO
IuoD2MVwmktNlj06OTYCwf2/W7oeHNPUa5umQOI0H+/C6whBn7Buxij9t6eq2+7Cn8Rd/BA54MZb
dgxEpqN79XJMS/lIsshLxp77qFd0wfXOX4rXV4WY6FcZTsdDZ5DkLA42kUVpUGCF03qxFu6E0Es6
UezxKSEAvEyxOZCN04ZqPY8X/uhDE/sNZmVHJ7k7H9LkVIo2uqH6WckqSH0fKypge+eOw904B3mA
QDgHY4LTQn866PaoPjzX9uwFAbfisfhD6+UdgXqFa3CkYyVBDeLvA9+SEN9vQePPFvZyDeeDyM/G
Fga9xqAehhD7lW461iIHUPZqex/aE9TdVEQIhQDX5piyWEBSBW2y0KxZ+bfGV+oKBA6kqxgzkLe9
FYZPpEWdXOVlEw5S/OgPk82CO0I7hg9tBScPru73Btz/zZXDrHRIegkKYA1EZ/dckZ+isIzVwE3s
uCogeBB2pNsoNK7uh4Vc2xH9djQdggyu1oEVvuMR3Yx/Gbr5GzHetYME/BZLMiPCbIc0AohjZzHp
eAqEH0fx/Ym40BCd/vMa86MdB7OJ3D6W7JCzli0dPBF3bVxfhmckGUiARYdpi10N+FZFpiF73IR9
nszniPveWwHdo2QYfynI3Ql8n6eKZHroJWOLjv4WsVhxQIlV024WpwvjLlorfdS1IQIvxgYqIeRJ
ejPvuU6j50//cQDOSdI6qSv+2WIj4eZ5jrnLf2db6DnBrhtZHLElmC4S2nKm8GU5FiV1HuzqtRjX
bsSpfjxbnchkGZd/wkeivSCmES43TP/hP8UD4dVgqErGjAstBdvZtCv7x5Z8S2VsUlBrYUEVbYqy
gcLQjav+vp2LLn8XQz0MtsFcH2BWGQB4ej+90CWu/43GqkpJ+EgeAeKoEqjju7oCBKgK5RPJceY3
Y8FeRifRoCJmb9WyhZ0UI/T3hWIFsDAT+V5ox0yDEX358vRaUtdPxR52/BjzgY5s3A0hzWTP8oG5
l86/qluY/r55KlywJenmgzCZXJKf1vFa1k8lxLsqy9bKyk7q48f5XpOUuNoeVepK6g4/rCV+IM/p
mg+maNA1CI628ZHba5atuLpItr19ZIeWyy0z2kRBLmpNiYLpq2moFkHJUHa0ejDPOf0jQWnOgvOn
v1V8yTlwpPHm3VVhkJ/5xKFbnub9bXhqVCMRyvmHGOo+NEVQuZ/Hv+OJpNRC4mlpz4JQWSfEkkOb
G/ozucpKpop3+cBYY5jM1KNScc4K1BQRW/5mUvCe+ElKvufTRZrwpIMSzrOHx9q8cJjyJePFmJeZ
RmkeKqdH+PP1N/mJR4+3p7EpQROOnf87zMr0FRJL0vaFFMGd410M1wpJY6M5dlKQMrYRyidnNqtF
LxsYQ7G2Rp2Mc2yJ4QmIHLCIcowzZQwyKKfjysuaOR8La2WNost6UVPW289CW1LmJuAu5SHX8Hlb
+HwujI2RjCaas4hW9CIlX7tw0TMCNKusYghuBbFw32QOHYmxyVCh7SS5MUTXui1pQ/tSj5Y9EFeB
WDsbJ8yQdr4FvhaVBCPtXXdsTfw1tJK8IDZuZ7Zp54a3Gvb6XakRaBDiOfF6+gNTmte/g48GYoPf
YSkwu77hlfwEFijvFvv6+rYMLKmqdXU2OlfrwTcMnoU63bEPJKn5O0c1PhYdCZfYFHff3aBwVhTe
NlGtWAPxNevK3osrDb+aZzZjhST8UWry5xBV3x46s7/m3GH/zTZprW/Z3icJpNc5bglTpeY6xO4y
lhDI0Gn55KIlFc9qMdqiv793WtQXYhNO/r7vbbgsPlZW4qBso9Ep47SQQQav4PPMZ0eadgmw0Q5L
jwSlNNTaurnSUz6BcLjLPEYJuDXitFhiXrO0Xn3tliWjZNH2ko/8y4Uj6+LR86i9yEKHAedv+Xyy
3X29Y1ZXOoTpN3HXdfa2CCGnngR0U6KRJlPJfiCK2OwemkAtTY+1EXQ5/n5jO7hXKU8ewjYevFUv
WUrNItaPuDS+G0s+A9yBIyNJlqfhKri+q634nnLgeTBO+fCXUrcyUwucPlQe24Pk9vXUQ7xXcZhE
Moru68a0a51uWYaimzHTlLs36UKbKYP95Ghd5q6tC51vmMdHWuFb9IuIOWCcv1L171whI1ZxCWuO
CxYMdJnN/uIEybptyMzzJyzxPDctbG2CUW84dSjV1PMNW22sy1Cu7xagAQxR1aEiOW9r3RxJ0uWQ
QjSLHx/eNltYmwVUk2SlVP58oSxXOVvVzAeE/QLPYlNkubaljjry9zTrtDjSV7J4HCYT8MdYr8sF
8GnThuFXppVzb7UCXUTpS9/ljwFq8bBXL1d96NExpl4Tkyh7jnszHmagArYWo2nTGSsHf3LFRLX2
MyOu22GraMLBNK+Fagj5wpHp9t9KTO5ccMoUjnYPV3fzzF6JbZqBS49nkOF4WiIDlLVHFuBvzTbx
qSBkKvVaadzG2gOxeL7kfn6lOyPJRuahNY5fIWLqMhExZIxIK5gRxrJ8Nsz5Uj+nk/LfWPugqiYj
OT46eCPOxBpkumyMR+I97aRcs1dhpN5e68Qge+xnj9g3mY0ko17dGLBvrAQBUDW609hff0LZwoM9
pn+JG3M9DXor/LMxjHAdo2olpJeg6wjiisEHPDLMmjQF0/TlqQc/iTbtqXol1eIbaags79UrUDPx
KQGUNjRkZNwgbOwgKIynr0vxOkDjCTDorrHfd53BrUSCDKkhiqsUcVhAbbuhnM/56Bo921HZmW39
WPKxE38fTNLF6OYX2mBl6NdpXh9uHvmzQY/SIXOWq3ddg3tSCEIjmRSR1nTCZkGM0ecXs715kgiY
GukidYsYyq9BsZu4AaHAPc6/9icZIB7PiKrsVZKSTW045vdmYbEYG3800t238RbQyt3ayVU5XTaF
9PR2A5zSqqyfChLD+wQY6oJaYJ/W5t62fw0A03SSUobH9V3oar7gSGSydMD+XyAgjarxXedSmW6Z
VbCF3BTuv6mrS5ppnN6/60ly5bJQTVCYE3KHZV6Eig2MKrQPtiJDD1FvBLa5QKFTM6aNuI2wQVw4
CXiTfGO4oaekrRxYYXdKux5UaZ8uLwFYAAX+Hg11wNoA/db9XFq9HAF/9HXpxa7xnsou90FxM/+/
4NHjbEGsArIJpdbvovodaC8xAVo0zALyGFK92Rig6y/NdXxR7Ha6ohv32DBfEPoPdrX3rPNqIpYH
Tq/pQ/do1NW9K1Bq027LEb14lp6kovH7KsDmdpeHRXIPBwQggQ11VcvlfpkLPsWTg0KvHUwywBlq
Hag1bq7qdR2OPfa8Yb1WyTIvtTNayGNJQZsFDE5nvww6tvYoSK8aoLeP7DUsfmJpGA/7xIpbIYW4
yubkRctXY42yrb71J3B+wcBhv7lRBnJ8UQRzolRDcJNW/F4dG4QnrZLCN3uRG+xRVHVRvnPjeveQ
OADnmK1aQ+pqgEzIl4qIi79Ho65pZ9+HsX3R4f+0rwFgB5JcdWNDjdqRN7aLOGnQt/q+MZrHHU8J
GBZ3sO7DUt822lPGdnGuIyIxechxLQh+EczxOQC4LLLQWQFmfHqqE74pKIDdfViInCwMuDga8alv
Dreww7SB/NJrB1inMGVqVAaVakpAzHRNzG+AeyG63dbqYfjqLkkAEHV6Cb2g5+9HoD5AqKofBcAO
t7ROHs7QSES7vXO3oSnpMq37dFevfa0HVdMJfU0vIrf/oGn5XxTonaDLZBNB9Wo1QKfYx+9FN61S
p3BWzQgoxkkbx8BuhWMJQNvCnkFIOBAkybCfx3Hm4uakCYg/w/Pb3SuEOtq+2PO5HyZEfGCew/me
ccgTvmbi/TVQdQT4G2qDBYeSEY/5utAUIIR+ValuYNLFuTP588jrMagIAhdTbPNyIHFmMyGboS+b
WhtiKH1Wpb3RQE0f2gCUkxn/ZP+ZgSkasqKIxY0Zql8o1XABYsirvr0Lg11hXzLKVvZEv8Jp2jfu
iKfFasUR5fmhLjS27O5f0RbZ/6tk4ug1h3Uh/elG41Ewy/2C0tZWVswwh3v7RR4T6QijQqR+XXH5
lSNBEQLE+/scnT8axAIdhaX05EarKJuydYcsHEAHb9okB/MBGyt8N1itqvOEv5IFDGTml+ZmfTUU
2EXwQchKiCfKlJb4PMmnjatdYyeur7EnNQXRXsFVMHXEN0Fosh2ONZeDcSVIgH9b1MlD2PY3B+gK
K9oIVTuArSczQ1XmWvdJRzE5H2ikZADpwdNSE1gT3ZtlsE+vXFm/bX6pZwPUZLyj8GgYkeOzx0/N
2bv3OnPRUhjB3drSqubAuYSVfvrQv08Lzo6FoSbIsLaRMT0nVb2pR9XcbbzkfhLBANUIpKEdHbJd
d7gwf5koDEYD4WAm5bb9RJdz09qtRAu405HnskG8/nKVt2hBT1Aav3W+YtnhVVNJnQikN77lgz31
xJGHPXbv5C0foY8XZpg0xa4yN5a5hwVJv4+xyU8MQhaH37xDJIrsRSzEXohkGYoBXhbp1Zweykny
+aLEw8ZgkKY3bsb/j1lYnmfagMzS8V2YPHWVnJgQmxqk6n/dooTn/LoO0OA+TSHogG32DJlMPWam
lsI9vRxx6ym5QGX/r9HcMPQ8S1bREN0YQUryqBNbVWgWOkdhYEQPMTk8+hdesTbi4wwuqXbY5Se0
qcsG8zU2XmZYoB0RDmoeTRJ+/3+MtBo2ewsQNyjrWrB6CbbxqBBA9bZevUmcZltGWSEOuwv+QQQW
g3klc0bBkOZhE8rj/hoBEKiFaGe9qFJYEOqZWDYiODzfAYzDe2SRGdKpPVK89OxNrkRfanRgpvgw
KoX0i2HYH7ekGC3sSSCgG+Unx0kjeEBfubSPcRpO2ek24Kf/r/wTN99622ZFfU6ORBzzDcwHLFle
0Uhl1ZgqMKSOSDXMbea3CF7zIpv1R2ABXvDdqQQs5tKVFLycdpUpcHFcvblKG+BRjxe0DLTD9P9A
ozyqZkZqhxFpy1Buc6AeGFQn36sgMrsmdYjRTQUZjUhrbnnNyiLIUn3EALPlU0inOY8dlxPVr/rt
yTJKZjs2xO0lJQbOu9U7cuackss/DkgT46HRc72l85sD5nbdazBySH78FaPKi0gUQ4OIItFvfWiR
EHUmdBMifr4WHVJQtDC8GH/xnlxrxr+GfTklAkS5SH7tf68AFDRcTeKCEmKUEPuE++r2qfzrNTpx
TRy+FA1a+XdEmaT5vyJvzqKn1dEFntELU+JcTTwIiO0mImrw458iA3xm8gu3kTozu5twRjrhr2Ku
ZEpdfdp529MbGOsjqTTuGSyNhYMZHQ9i45nwRLazZBq7jEEPUPVsb/kz6RTFTeKzc3Z1LuEkJnIX
Ec6MhhcsD5R8w3qMfkgwMVagn19qo3oRb29TrpggMzvH2k4xLhQvRKxUS7LuwMjQqkJsj9Xk4rqG
DQt4di3Ku5fuhcOKFNI+IYcY6/MXgIij3flRvdc8b1FuKXSaJLIHBk5kgLy3n3kV+VWgYbBmNzdv
mw3F5+R2HwF2iZA/P6o4SxadH49JtgtkvqFzWafF/2hz9dt9wTFGByu4CKySjwOpNqaiRMtIcmm0
hvorr64k8cNO6s8bCFNaZEtODsOfQshqbx+YsRgT34G3X1EF0PXNvJD9vRnwBZw6uJqiUDRyYg1r
ry0CUNYIpAj6zPfBEPQGGaFdDkUX9vOam13VDuKJqNl9z79Wwu3pOcYXMcDy9USpf9sel2Zj7SkS
4uRDYr0vT6dWTwM9/bX+dKdczjxDaMZtXZD8dzzcmDnPQDKDVqVpNjXa3zJscBrpw3s4ftlNBWJF
2LwzwLU+FTsiGWWvJIUdArOfdujVsQNT6dxhLd6I1GE5FevCymuIBhKlPvJ6No/vj0MGCDA7+bit
XsdPyAj9Q+MLc2eVjI8wNXEVg+BX6eQZh443Rvtpb98BmFjx0Dr3XpT3FI27vCEU0647kdIblA/9
VEG+ghl6kYVdnsgKdUV7aYb5u6Q+18ZuQA1/3VfD2vXVYUQjxTtKddW2kIHAwF/Vca4L7G1Hlvw9
hWMk3JLmN/dkI8rivE8gYaBQGzv8zsejkTwhWErUX1lPfoMvCZmlyzCB5aPt//eDI8eqorqzbYkS
hNhF+TGBP8iG9QuxgNJeZBNKeJbbJbBB9CJRINEqFD9h0X3cI9yb8iM3p9og4zwbZ8C24rXzAWNp
eILj6mGi0vbOgXfrhlSuB67YodV8Hv0Hp17FZMXNQBjlazqVMaiLfqveFB2G0wQmtdlvpwEzqQ7q
YgH0ZgjPqoXFpukEUa5QsJst7IU1zFuzAQLRJeku5n4GtlwSp4JFjoI6e9388B438kn2xX51+nFt
URWLwwUI4gmDFmoDyTiGj182sXTD3qtJ/i07wQpC4ns+wYoscFEZOlQcf1ag4XHv3sB9rxbKVOpK
mcgsA8vjLfFlMaBNd9eGKyf9vxEw1c7sUKEPvSGXvXusGhlewvHw9R2rpqQ9m0uDwPp/Ye/L6x8D
drPVIpVWt9+eEUAIeutu3yf5d1mymKNRJV4HND4C3wIRyZpS4dPA+VP107trRIFgDiu/A3cWWtC7
/mkP4euLHHjKb4r02ZJOE5Cs9vvEnBga26VBMRm94SBGlFYyNQLW14OyF8Y0r+3UQL3LVNtRgMmU
VGRires0GG6+bVoR3THQil9Ixj09SYbYLWk5SicNjEn/OeTHVheL4r8qjW/2y7XEmjX4/q/96Q8y
F4GwQoHmDWefUeeAGy5+/Kl+LAtIGspyvwuKyhuKU6C0ly7Bu/O58JpGvPH2XuzSz0THshRMphCg
zcu5ikdtyJeuWeZ1jU8/Z46Uhf4QBDEul1AZkW/LJ3yDhA11eH2FJlZcQ6IE3x0yQAycrLYdqiEB
J5u/aE4HnhIzkqkXv+fkzdoXzPNlAMjzCFLhN50QDkwlEfShbQ/LL3taVk0xjpIF5kwm70ghbOV8
+KPigg4pX6JrH8Dhjdr7Z3mAHVuuvEDOIoQulXWyWp0nd34SR8b5tLJ7leUPAdPzFQPnchOW+UDo
1BANRfMRvhESHz4Sa4W8ttdOD/5SKC5pphEjRFevd3ohoQaIW4XhApqosRD39vRu7sITODNiCqEz
33jWuPNJ7lsH0uzA360UjzNFspjjFggC7l+PXh3Y+qM8TZ9JZD2GBYFxvYN6kpk9Jq5CdjeGIUki
qicfyITIjr8hxhqKwoxKniM6D/CUB7x1sUQVrorCF1jD3eqhCvU+zKab+IFdUW/aCN4YhgP672pd
jB+C+VpR2KfvH5TZkdiiY7PNZHoQwxKopiLkLq46DZvcYIk5Uy4NhjglYgwTwfKeZv1ehpGD9Bqi
5BVZeiM9dEFb8Laaqm31UHmJ1QnUcYjouBnMk1rKv90MISpPjX9CaFpjORgRDJneTwmqr4e9oOZZ
3xOuSbpfI8xR178L+0HmOeu2HbXrgJzz4/4txHL6OGftlUGyBurgyAj82qPI8CLpno7Ik/paMelF
Rj5WffchybeeG1dgwORvkTqRlFh/wIbkC/LUDbaVa4KyuhSQiiIP2lMtddJ6Dql8ReBN3f6cyWxC
pNQz+xcukvQFQq34+Zy4PUwruzl+OnRW3jo8Tn6qqc+r9+TCkXnctDf1hSPnBQolrPpgQDdpx9fZ
mEc1xB4Q9p7niyLoKOSOuiE4+Sf3XsV5lp4+ac8FE8e9uleZqjB3/sn2lcYK502P8EFZZoSgVz7S
8Tk2c8hrk4ozbXqEk3/HWbvH4/FE5GSHl9/8p1aePeQQx/69SQlKG95XiyE3MBMBX89N9JImjsZf
kJ7ZNK/k99D9rDCEzbvzejCF3J9FcIQPEi7C54vME1bOYPShxvybkRIatTTYpDan2h9qYgC7N21L
MwKhL1sLN3+QtntR6fAFiY+A+c4Ht+qHvciYPADMwdUgUw8mN0+ZwWSbd4fJCXkAFaYIx8qNKwfC
Fnh/2vpCpyN8y5FPYTgdpfNgLE7AF1uOaHBMAP0dWb5zH/ATSEORwj2cJeMMA1PaPHqLSY8qfN+9
mhKsvmq35HE0+21oRudwtczQfvnYR5fdImMo2/T2tkO6SQYc7ZZ1urWVXs2ecGG/pAGxJWBXk9XB
Lg6gy53k8ZGZ29433c5rPOIBIjEar++Jc/Je/G41MqDnBRQ4MylVkUMqlRo36wMo9Z0znfeziov/
id/dMVc4Eb9wUqS8eju6oHh6NsMdLIL8mMpdMGZ8ffjReTqO/r+Nm8yhub0Yw98TSPphIq6Oq8lC
Bqmuq8q7CKe3MRde3OGavND5vgejE4K7aBR1DwI0KafwHvX7SwKO9qyE7mqBpkB0NdYIhK5O9l0X
rxzKALnYwlhaiNDiBTGIohZSWiGUDvXjDF5ehh+KfzXUuVXPaaBtuTu5ZKbzQLbTYb/irvj03D6Z
tHoXTZTfhWkCat2Fv0FzqQusQZOOjPyQhmHnusoLlqD0/qSfPMNXJCv8L8ljX6KQutC02UER3Iaj
RTQQuZv+nMbERZ4g6kjycbXJ5dZCdS6y5PSB2ERhppkdXwkQHbUbISOhOgJpOsPZzT9qZm12knsj
LJtPui+DbBJhxEnGAMjr+G/xwEDxdFovC6QKbbYxIKC8SfWLt6/edIiwjro9ZlMlMPHSuOAXmx5S
Biz/uXMvJLnQITSUTPuloUAB3iliApB75MJWbxWejQ8zcWyaUp65J6ceUTp/8Og1S8qnDblQFYAh
uTFW9J4mXyo+2fsB/aEDwjMqmh6kpK7uVIu+5mK8Nedkw/r6JpGHNFRN2xpgbaU71MdRR+vRsuaK
ZjuLEQIo1y8ucjFfoxXct9iJPXYqNn92SKlG8Zzfz+23xK/cw/Fl7UsELz31RUWowGNnNirjXFqz
/lQQBGfjiAgHQHJBc3RmDzWk32WRHwoNhqpmv1I3MZ7B41HAKRmy5guBv7PH4oUfd1dwVgJ5w6k5
3ze8OgQznFsKILxnz/9uWHAVskhQIZrnbHl0oNyPD5OtGz/Tu0hOU4TPGH8U8qpV5LFBCsws7UBF
Hxq3/ZvM46aIoz0yLtWhv5DCyV8J5nLCw/CiwyyrBjUnyoRrw32g0rAxFf7d87/eYK4L3fSNc9Qn
gClzTxJeSnwynqtLPzhv29nuzPSm9NfdIaV1fTiZM9xLOXLVUBLCMUxq7lOzPq9pPKepjRg+izys
HWwemMqlBK0/njPRtBLaHlvYjuGHb0UT/Jkq1/4KlfIfE/s5HdSKLnd3yYYB8GISuHNDtOeZRsiR
psH/BA1wymI7rZ32YoFU94I/jMn1d58evfg34Pg9K3pqy4amd7xDSYntqMujrab+Q//746Ry1Yk8
BCR0VFlg3imrMtlHi8EbUF0SRaC0tlWhaQ/FWC5BxyGIhnGDiOBxqE/HqUCv+7cyoQoY4rolAdEA
Ec2LHeVZQPMlznWV31tjctSMm9cOL5JwnvS7/ZpEHZeN4HhuB2RdMSsR3EV01DM6bTU4AYD2Vmvu
NdE4PA4FFlbWlazfmS/+h09kchXz8JtN6W7jx9zBYlVZ2HXxfMU2cVlfxhgCI451hiH95z6e8bxs
pI1Ivx4BqmpJ7g9wIQxQS+4srwd9kRDN127rOSd6HU3TdjQJIGtDeoHrks/cpsh9EplnMebsq9zy
gNET0YI/WlRKdk7bDU87oUSts7I2uyeWTngFUrnsdtqg1kJSsZZCH2ICT9VeyRPBZiokuOkPmwmJ
txPqoZRNkj/0p06/P3EqiqEi2NpHipCr6876qAVe+LnoI5n8VUHiYqVYiQv0rCEhinA/avRUfwbb
eos7NfI46i4UMWH+jKmYdDdeae3vnvuesWjsIhYqhi4vTeDMBZW1dwxIPCULhOH7vS07jG0icEoK
wm8NWIvcbVK2/TI5mHB5EvOPr53P+u3P4LQv7bVawJr43hf63WBjiWHVdn6rWoMndYwqIyVQfdVL
9TpUWPZAX3upo3gdawoR/74JLHA7FHluUN0oK7tPTmiMjuKiw+I99mHLRX5fHi4OP/IXRoDDMWMl
uy5/2JPyPaIshxTe2O6N5ZmzL+Q+iW3jckKR03AYNkHkTwwrmkpEKliUc3wug+WyBJpsqCubEaA2
QPZX/E/08Z9iH1CiLvf8PQQi1J+lMb7ZytKdsYp3ZgxQWkz0DXreGiDNeFlmLs/eyjYCjYOS7J1d
iMwTu7J4MZRtQLvJ8zj2gFBgs+dW7njvJa58CadJfoRTM8L86NT36NVUPq3qC7cw9ntjWbJzenK6
sNPgZJGLqMPxovhn/43Ai7Evj1yQg4LXxs2/4N8Yq8nkZxO+P+EDV6/Q98AvaJwBdlTHtoVd1E/s
ODl2OLKXq++7lpFr7lJIwR85bjFZBtIt6Qo3wssXGutmhphu5uWBSxK1FCsbHOpb4FztTdlfIR7R
hU+04jkot5knKlOovlajbd0wpwY3O3LjthtPkxwKr8tXMG7nBgKF6xVemnaa+ZSIOqFlEMLh+Wyk
xBtWFfjUmTt6TW+nVoBbZXM+VP/WZZgHu+ccNJYLbbSmeJ4oyATC3gbKqY6sJi6hevn2ZGRc9K9x
KPomOhccxk2kBr/1nvHFNeWqBeKNU9n5I6Ck29kh2dGCM3YteS4DwzN/Xo1dTvZoM+JrpHzJkwt7
4Fsr42omBtg51akjm8aM7ebf+PcaY125Vx/myPLqCoREikQvycQsiszOGXJt6KYcBGGgV+FrFwgL
TyCRQeZ3OU2oVWkhGgJeqZYqnYdAU+Wipd3L4RtLxPhOoxpW0yJ20ZvXK01PK2h+u+OycCJxWbx/
0AaXnqllhLYFGoQhD8uhjB5D8c65xfnu+ySM5dDFjTsl7TfIcYyYgZqpg/3OTVrwO/zJAt8I26El
s+oWZ2yubcrNV0SQ4wEWo6l55kljKz6ztwVrSjDV2E9YYV69dloLcKEiQ6/kKzKAL9wGhZleVkC7
6/M81V/8JIeTIcSuNLBslUOmeN+TMU1UrrUR1s6N7v2Zqg+cg2S+FpcfSMxTQnYXYeH1wEpwrXx8
DmA8tg8GTr/f/uC/f+sUoDptZRKX8PqDm1kw4bBVhrVDu6ASgbbw0HygIZ4lECeXRnRCHXs9+7uh
iocJGWb0CUzbMgr3Zl5zPlCXVFMR/AlT8JX/kZ4CmLmhOb7AohCBUqDTLPMovZAvdrUmsSgQDkxu
DfyupPPh1nEVID6xVARaPFXxtpp7JJiNnUX610XX8XQQc1GwaDDfoAEBnw40f95vdP/SkxtcPre3
EtqUQNXamL0mP4zXi8kNxehq2xlcniJ0UrgmtOQb58QwY3lRI1yI7As0h7KkyNU8HjkD+sBoD70t
r9V8DF6GkkZjCeoDJEm1PRQ7oqNJy1bBp/Sa5pgZqhD0Ha/Mx/aXxcgk49g/tDaqyTAbFRnYw8YO
lyCLdNVgUAr3G/DoRxIKJz1I37g6R6CotLUGJ8lrRCux9n8l6+hJFAWOz+IcmqJvuLAnnguPOYqh
ElS5Hj5M4qNwOFBHO2QqBS7MdBQScZDL6HOJOgJdBLiPYwsClaKscq5Yu/LTrPBlDP2tcXe175wr
jtTkQllADOGGoWbepyzAwc5ahemapzRpQq3nIMnSZFatIDRP+OAL4AOsylWF6oOTzJ6WO0eUiVQk
qwRU1F4mq+HvlfzMGgrm24eoL9eHUnSvOE0387IFZSfnmhFKYVYn4KHMRcABUCtdB1D1jHWA/1ix
orMOnUHzb6XG0Xr/Y292HbTiYPSlbP4ZE8mYKRk4wCweGhG5HDnVKOpgM7ydX+roSzbHfzymbWw9
LLdq5t6BpPcFBkYx4Hu+unrOD2ooKaJ7Quauy/Jfs/SJmBvF3UaNNWSrjWi82jP14/9/F9zrSiNd
RANDMEa/qFnVpM26i6nhAnBsZA+3t+DQmsnl2QUGHSJZG/TMm5n8N2YD0P/qPuY8xPO6OrmNUq69
VDa5wg5cRHRBEs2l6Nw0jCHANWKtDybZtdaQjztSOZlRMue6MwakStrVCJMRuWNMjVqMm3Qbc5uG
GsrKq5/fy/j9ODNsWApG/0lzJmUH3a3l4XQ4vaAfZI1OFL5a85+NfE8qzgaDoKyWmm/cIfJGOD7r
Q32zhyWNISPL3tqJgXTJihB2qws8ig1/PmBt65Lrgo9r6W45DK0w73ASQk7oUkLDZZNYxzuyg/9F
POhZimWdBA78cx3/jfvcDYCOYyXHofejSV8x3IbHAmtuZX/m3VhySde0Sg1EcQKCwqlzp71cXD6T
keNk7h3XHnjdBHARoOp4PeUsRrdxtvrJsoS0Fj92nQyY36Sa+r6AtJml+f6aOOQAIqLOhc8xTDZ5
tqNaSuTZtIVlhNMigOIwt/xQ7xzbsnBSm6wZJb04TRIWO9N0WL0N/0jOW9xVrTK54e9bRnJ/0LDJ
F+Jz9euxBITiaXnJaGczRNnJs+f2RboUfVtgfSCS9N4AvhQf+HUp+B8s9NLf40HS0qzOtZvFfmsO
a6djCNpGXX9VKA2UcVJxcSBFisTouiXY3235a0M3Z0BD6FUvi5BYCU4LNDzCqhslzJu47/PH/C3c
oR19E19oZqGcI0DIsKt1sbtypids8YhtQWsKx7deF9KDh2T9EpuIe1S/bjBp31P9Pm7IPdah7lio
o6muCC81LwX4tXkxHNCCswdDUWt5CkTysCFQTjQy2lLP3zPrEGiQ2ZSrXGm2uWRLcNfOEk8D53I5
Y2wXlEyFsVIe5n+YoLV8RKkSyYWWuDLfFs6zLmjM21dJziWF1uyEjF/9yRDY4cpdtvFk2BPVe35E
3qIHGFISdsh472dtouop97QCHD7WcWp0Z0UnAvHrto0v+bBuJSrcHzOKclw0reXOBWkahFMft58i
AH+ZLQsJXHTTbf32myRHo3d4l9M9bKlJHlmRBsW+2HyUjqJUgqQo+YAw2P4zrdt78aHxlDkJMo2O
xcS3VPZ2s1S1V8Zh9EObOnt1D66atWoslsfK1OsR7k16O3C+9E8NhnfeGElVvGwtHNf35mcNt22g
IX3ZSN9X3tNG8Ri7Rb4W2MqDzi7W/+WkLLNSp7KK10UuDt9cMs2QgicpimDiOsKXDBUS4x2o+kAe
IxyVY6YvibCqhsLKbH1M5tV+jMUrWyVRRzPRmys9bkwEdXitS9C9kPXCgJHQxG90quNnRArtCuS7
kdjTMQ6sgz+v2B7L/oI6fEnFZmdGuxfeHWcpJVDNpIOVz0dedpCD4YlHIYmYgNspU3VYML82lXgQ
glESu1AzUvKQlSBsaSNV2D9wZFmDPUSXeutXBqdoZlBqW153uLYleMvRk1om3KRVw3MRl++3rwVz
hmFerWJZUNNDR7nY/M/lGqvUIe5qCDC5cLsFLlNTk936wwkyqRg6GIWTjJXl6vTldH8/EVI1UPkz
GF03BqwZtnYdgUmncfzO/QIX9nQz3DQCKDKFXFBuZh2P7AgHOaew70u/51X+cBznzkfzeEoqRNNl
DMsVXTaQ6hjvbmXbhLah+JmNGnieVSXZwwYPSA+uWuq2wg+73TgB3Q7DYtwn6wH2HEaH+m7Q3LO3
r7TJ6vb+Z17HzYJdENlbBsZSbgVZBgP9JbAFLKG3Dj7p4t0Lr9r7LBTImKfBrxQnvpiwqd7lJGaN
9DH2rkS8aAL4ZQx5xPcSjmjz1S6VeizPOQCRZ1V3tkC4MY52ZmSeNTTCIyPyIR0h8Kam38QZqhE3
2Zom4BLOTjwjCRf9zO5a4lt5NVVBL/4yGcjYMkD6DR471m/fwxUfnpnbJuRBEzP9Ypomy7zzUzp4
0ycYwdowG30WOZjul8ZPZl0Xu9GU8EllgD2dLBVRU3rytBmQ7iD4rmz8ISxYw7zSfArp+RfbcRsO
9JaoRBiIIxJVr5Bo4MtE7V6vaAAqpciDkrDnNHCq1l7X1yUSHx8yc1zScsL0il+Jv2qPS3lg6Sjx
soiczs14UD6I50/2SC67iebNIZpJ+iDDCfyWEg/ZOGZy+ZSEtj+w5uZGhDM5FG2yrB+WkbstdmH7
cvpark7tPPTpIF+FSvYTzfHzj+V+7nnmQFQMf4tqZ23b9ML/284wGHXFnMGywpNGquYbqpwXLNCx
/AbPes62nPBomgnbUuHC0L4fk/8M0IiyiuhYl9iX4izon7R4cjtyFdFK29Gc4W6Sis2sKbnbsSMH
QwkA5jQP4IytUjp3y8vylTbL16FtKyV0su2Z10ZsY3uzaijMfh0/2obNZLpxFuNgwGrTNZd2El1N
w2mchA5jlvG36RNOa3gVTmlBM6zC4XTRrg/DAjIaNzhCgMTEx+HkYi+23aWUvnjcPUP5qyeQP0Rc
G+2PGezYBocm5UyUQ+W6hVpDVqEQiVMM9v2URWtO2oFmoFadVNM0JOMHwWbdhWI37GPCDnAPOtbC
ELU0/mRIBfZheznnLgsqRbIxM4gvZQgQpEtGlum6RZl3wfW/jO9i1TdpMVnC+k25ki4lJltjCGUg
BDfNhgMDdnRbBPXA1J1DSIHVfFJq5RpsMmKgmpU5fheHVxdOROwrW9XcnerSC+49LIg9ohkMIvZ1
MczBgscyXyYuANMiUUwg2WcNCkUYA0E1oZiAAvxCV6E9xiK3Z6pMGtVXWZgs+TnlApE7DOkPkq0M
VWIeS3CQtPyPztc2pxdacWcTd34PPcQR8WTu69cSl4YLV03PepvFcqX3LJmByUCMX5Gi855Wu33c
CaX18a8W+JdTkH/dpg5rY+t+KptdcX2gBXdjGhnlGbX3QqoPWV4XRNPBc6TjKuojHvGIMz8dap48
RxtCAV64YexOUJaYu3lc/KPr+S+PaDfK9FkCC9NSLX1xF1IVV6/kfNGbmZEeMzoZ2aQVs/m32bcy
iMiUwPupZNf1HdPbPsrO30PSSX71jASMT9/qTmEA5ZDu7fTRnCyV24CnPXPIrhulbzdyN8WzWiTY
c6su89t7r0dA8H+aQafj50MUr6xN1CZp4/Pyfqmon4fP+ZFPh5Ynb7JD9yOO3nM89qaubVKsdIXm
LhzHXY6FQ7N9jXBdNwZ0Cqc3InnEiopfBm+JPoUmDNSpQuUQRdotFc1DmRTBrRzHeynhItMV/kqy
bGld44l3M0ts+0MYsydcsuZtdGuYu5cilXRsn1i5lgNWzGidkZ/edRWq9AKCtSQ1GwCrfKahMEJe
EN5tAYKQIHm5lBR8i1koLFO9XCZzuSDCxE9AvKjbZo9UQTMuOCVLCJCR64bbyF3os9xCu1WV8Nw1
1xnwLMC+C8tZyr6zaMmAI12tgZkTsyiwQBElLyYRLneoD6Hh2Mtiep/NOcz07ebS1IgLpXtdI4Qo
8YCqcu+0JgiXqDkm4u4Mjg5EJZR3B3BtLjvuugBY/yl65T6pArfpeFwHRf0yOZb43CvL0Uw8DuLN
ZWRzQAPNazYTSSiDRFHDa9spKEjsMmdakvyIebesuI5npjGKehMZ5i4eeS6is22GQAsRoyTMJ9/L
ivXNNcVaTJDgWmjSobxKZzfjsoXLGLfPigI8yJWh6Cs9h46UQws1uvwcIiroaai29vU/ffZQXQDc
Zi/dq8gJg+cNV8IUX3cb//8FKOl/F3khwYK93MszOtPSoqd+0BazaRa17dzpPSFQJpurmFpADZyk
mchBj76NZ8Io/PKLQ+Gl0W0Vu1x4Fqmm5De4cBmhEsPqma86t3uHexzx5NnfccbxUYvyzNZBYEJv
YzY/7mu1zNIucVFd60PxRH5N0kLljs2PcIUhSDHYsCb4n46RuR0K5xwZoDzf/aH3cRDVOjZPQppM
DPsoV2cUeDkAWr1NUJ/WWe2fjUZI3nv/bCx94QErX8thVuVd8J0dpJ1WzRRyZ9Jix0mKGKdJoNoE
j+9ZHQivUPpg/V3xe0vyB9gHTL2ZA+6gxkXJiKXObxU8j2lRfYPt3fcxE58AERHQ1mDWSsHaoi4H
npXtmv56P+c+1DlNhWAs5mdl/y2wHKhCWJfYM2gYF4/6ZnSCYzy3Quc7Uaj/3zeAsG9jju3KypAm
dftiW4Aw5U7ecYSnp7ma1qwcM/VjbLSV0Y75fSaeZmzkAPD8cz+Yozxe1XAKYcbSjJUvOsdNubYV
61fNsArXXpO+dTaasjH4nW6gJJkD0zLR/1CteQ7DbukCfG21Dq1MR1cYbldXz8AiwD/Wg6bfIrul
Dz6BqAUMeEYoLj9cTvKHNJwOXrBScI24TI+ZoLfmU/uEV4ienUu9ibUHkCa0JGSQX5bLwzPcd6AP
uKaVWUYT8xovnBPq1RPNYMabHFWEE+PyJEqEWwv1V1RUa9BlpMKk5b1Sg/7vPGJuriSQuCHQsm4+
5RbBze6ud1eUljE4dKdd1ixm+mooiVj5LuJkr3RZzgh+vbb0OeCRS+LS02Cn4K0QMMLf8kb/EiSB
lqzh9bN6k65N1UjyOrN/skfYf5uexrmwHr0JNhz7ckNfSzi2jNAZE/0EdLx7x361tfqDKHlQF5fC
Ra1qAO1igP5YueEBGA0S1Tz24Icez9ew39n+KAHdMtd2WTwGs0VnigjunAx/rJZE7BvvXGC+BtvG
YXKqLrpmYmOmLc+vjRT43P7+dWKn8fmW+irLailoGDmbhIvfzraFdCRZBncoA9zISZmQUqT6lm+u
kK5bICjhw8fgrv2KPkKPqI7iKDg8NHio16zcqEqatPfxiiEPikQtSS4u/LfUBVeYvE7g6bUIOQd7
Jm/cuXVk/5N9BzDzYRQvN+ehL2QNMRFVNiqO8ztFweWspORSf2oEm95W8JDOg3T6fnVJEtFQer78
DPdKlC9GFqF9sp1zEsMNqkqEcgyTzqvyV8OOoo0MilP8pAexJqk3a5ye1yrq3JgPpZfgnMFSzJfF
kWEMhJzij7EGkqgPW0VcW+MxKE2wuvNk7n+NIht3i8iOT5IQrqOwQFxuDx9MTUIdS3/a0cvy1KwE
gUc+1bCLCmamKBVPsLT/g4QdKTed6UfAnF/S438wWMYPDokoWXCzl8wrUZXTe4LqHccHXPwI8uBt
rB4aIqnbNCIRdFvpQTxnoZywMZepZO1psCk0lw0WZ+dHo/76U1H+lS8I5LGPITYdaQZ2nR+zot5N
zSNiG6KGCjTgRbmVrsgpZL01jiVfh3beWqP95LiBQSW1JbPezAlr/QZEvIDzerkQCreldjo3muzD
ugMtLQzIyCBHmgRJ/+umXeLEIwGI6ttZ20Xjl0eIs1ULyXjKgzkj7MGuLuX95xxtbzPkHZqGhtH5
O2gFdC4W28LVZQ2coxVM/f3fyBQPm3sYE/5YXaG8NQsATQfq729wKKhn5hc41mkCe55bB62ar1w7
GGxGZyLjzcCBZSV0VYLNHy44CSOvUUKcw0oUNQNVQd7RiFcxIQmn9KACe/NxoaPegKNvSkrYRGJa
vXrLeGfiz3rrxc9akIxuxjbVIzQOdXRpN06Z9iYcGMYpu+mCQVxb8NbcORTpEm1cikVcVFAnMBqT
bjZWo10sZoOUH6E7iMkUp2Z5jremnyAFy1uuEuE76NCG9OuP+/aVFSTyOAtCk3+jb4TtVRPIKqHf
WhjiNISbVhBZr1V5ruC4Hnw98DdnI5YVwKv8wjUxaTwj9MmUz2E6DzQ8zA0xHBkrIFj7YdNKj7sU
KDc8AT+ZhnuvZYLLJW+brS9gS78UY+Q9jhmZvZ8/pXJK7N/KmOq4z77GaJDAxLlB2CmWJwcgvicl
y0LeoJzEJEjb9RpuD9pThN59enPcgyMe+na6SMt3DUvhC+2LbZLJ1DNkTGXTCHaxjEcprkfWhkVT
nWNB7TZwEMJsgCRUuEPNCu728Y154/OxeLwN7fWh0Ed7YR58DKF7BbjrEG87O0A+G3WeLcjjCIyw
rdrvZWMhU52OGTQQI9V+grJvICtz+51sEPjRgY2yNgec8/G7xHutSkGSTAfzKpQ6MSY+T2h9OZpf
k73VFh38qAjGK5ZZ6hZsxB2gwyqRtokLgCZh7xjzUMeqQbz/v2jx2a0H0qTXidzSV2tPqkcISHED
q0cgBPyjcqC/nKstZwpnEvwGUA6DhzVHtJIcguOAWknDC5jCiBifBnWdVfK6eQZYXsk23YBbLV9g
dMRqe2t1GENpPpQCaTz+un/GJ+ruCrQz2cDtAsCwDcQzJwkewYOmThat6NzbBos3Hzmlli8X9Htd
pFCHSJ8Eaw6QCfQ5aXhEnu5GR/tIToK+OS24T1p1YJk1EGTuX45dBiMbipViyPcQcc5EOzbTONZh
ojAT/h/CEOjJHZ/q6SZGzi9afW4gEZZSSiUmh6DPmjnhzEMv9XmpbsC/+FYhoPzKVAe+nQVFJ4zJ
L7n2+aMz2g4WPTT5Ikdz2uvVduOsOYfP5+xDPdwKNhSo6ga7N342woemwOmAPcgcD7UFlSle97TM
3yD7epvHFXftNTaEKKg70jcpqWX5xPEdagxOiznzKNEfq5ck+E91ERh4v/f3WnBLv+C6bXlK5rnK
bBOaEBfzcDf+X0qrQWX2dKTiq82QR6u85vnYbY1gh6n6WxrdATOd71KgSmFc4XO6toi9NmjkiNtD
8eC8JhjAXxMpSVpVGUpnFgKB9KCZTNN/HWBEUIYD7APotzBRg7ca+Oh3+WMMdJX3KAC2SaMDLZK9
nAOqI+7DZj7WBZctCCitDUn9gh5j7LFKmYyQf02yuxLBveQptbLXVuyhaeeVLGPjTI1yGccNVkCl
jugMdwzpuDz3IKiN+mVpFmWeUEuV+8qUIOuWbeW3tA8rzLpi+cVnsziNRkIxFfvMlEekOmmonM3g
0Uip9hxLGhjKTuKL45ld5e91xkQwwd4wjgHV5gedKyDTjKvCYy7THaJrvfQzmXg/GUNd0vePwoWn
BQp65n8OJ2EsDauodurS5GNru0FWvvekAG4UWIWgVXatGndxEE9XjWMJKaheHvHo4xhlsSETdZx/
mrfJy9aIgaSghiBaxs/S9rHKPBm2fm9vyg/Xs2aTSUk5J7EJfuaixEaWtfDpxXEhbI7pNsmDffu7
D1FUVcCw9kJztRMctF0KCoLhkIPXGyPgJ5SgcvvNV9K8SOi3q8HQ8BELsyVFdI9HTHZScZ7UK/Hz
pEu7YAZ6+7id5SkowRZ39DvPf6+A45Uu3rpt/FLcqcJ+tOrplPa+2v0hjYeGnUlytVo0+M+VJ5q+
zeTKyDs9NNr5l6EjdiUnxlNJkCb8NIVwmjrMTc0fSMpSc7e7rWdoDbJSTHAcQTRslv3CbiBxuUe3
VdnXRVU6VpeK6ux9Axp9m9w2Oh9wr4daC2oUnbeOjPHnNOI/x+P47MyGaQyDmqLkeT63wpXscWAh
W/NzLeoZK/V0+WjHopYE7OMFu67fkB5xF2IsaJ2D9pUmwU+LI221qi/p1QQTL1CftvnNmLa8wdNw
WAOADOcdDuTC6XLfjLTe4gYwowaPH5oWOFNl3AZixoRa+kcfnyfSD0rLZZmyGBTv+7zPYf9bL8+t
P2ENJ84fI14IJH4gmcmzljPKtbb1+vXo474CDGV6yibS8nVRZwVEVmQlywC3KUrk+H8EeRQomnlF
CYxEfUyU0kCAcdr431yh1CYU3bsrwqL78yCz66c2Lavl8cZRMn6XAeCYdOkrucLIzPIyl1dm7Uyv
9daBSuG8UnPoVwkKAMCCNbe3ox3GRVcDGcOhZr193ijB15i8qV82cv+j3TlbtI2cp4kTiwknvL1P
Bp/8+mff6KOEF7wXzooJVHBOJbRwXZqYgvZGxWYZqdpEE3IvXl6eZ1bStOagoFAWVqC/cKtGUESF
rvdu0fVYshfRVhnCoaZfUUnc6405NGw79x6JlcK7ghhG2mdN0dg3xSMMAl32nbOhTX68sOtHzbk0
d+EtidosKquPW8mHEYNkvHbZVcmgGWn5C2/PoBcLieq3vrgykgIEHiXpG2ciirKQ5Ngw33aXE0+o
BiJqSMg2gsOkSC4y7PF4c5qRiClRL5G/nDZm/mIRnwq+nOduE6X3UQp8+cZLZwPP45ygS5+WNbHm
ZDnxBEQN9A+MGu/9rS4NOQy3/BzEgHyF5DdJb6eqmAFS2ja0l+cHaUSTEUb8Z9rsFNhW4ZjnD4Mz
ZuSDVFFaLhHSY71mD05XZCdwU5oY2uwtqTg0mZ8o/jrrnMFS2O77IKm+Zg3ocylhgNY3Gj1VxTGU
9//gV4q2LDzMErkkZ2WthYCQJCeWqdlOfJSordoPjALicDNz814ncqNQaA/oyiXjhYC+6VFle2OZ
fPYyf3D0uxCKDj4PpclkPHVm+wini8ICRch8HbCqgxNeo7ViLMbGQJ8Q7wQS2YQEexacTq4qk+xS
VCG4Hokj8osfuEWRfqmcMRtyFa8jBKTlL1hh2op/Yf+r7m9aW7DZRqtyGPA+4dt/rnwFVOtNH3z/
onf7fo0s43qIXacQNwRiTiKiUeBxlendnotLT8jNCLFvuFH7vYdxMBaQCoFfTaiM2KgQZsi/OPgb
vk3fmJPfeIGLrHC5EOkBwtr1TOf/EoCi/Bl9s+dUvbQ/DECQf/SaucVDIzWiaG5HhKeuNKFkopWk
qrvmvDNXHqz5fbBHwKjcZ9rntSyvuyzrz30tJPQ6lrukh2NEAbHtZOZv5RyGOF+UhErbs8dcIrpQ
579ARJBdBGsbcgRb4RqF5pN5dqHMpaCqm/z8f8he8o2YQUlutYTycUmdXRgHOQjkH8IqJO3N8KDp
V+EagnfrZLlwhmaxoMkIQWfRwT01u0wAtB9oTylR7gEtEtpuTj97wW+5B5FgryjhG3MwmGpygsNo
Ex62jG1MPW7KRW39vmdAimcf1V9MPP2e8innjbwuYZDvRTG3kzkeYNmt5vM8WCySjJlUSS2wn7IW
v40PPFr58gK+9qt+yVNULSRPIiZkvhflgH96hN1nJo9NccgHlLOlQpWeUHUiSZ1NxzBinDLo7vef
6yd2JE67zjSaDhKSC0XV9sDI5HPqP8fzPbfeuBJGTU4dVcvIT54P1BK1nDwxT00/495SGqVc32qC
Hzvw5VDR2Aci8k9x3QRlI5ToE5X5c42enYE+ayvfEdtRSOtnGLidC4pJFkBIk4fhoWi1zyOICXIn
rPBIWsmMFJIUy/pKZJCQo6FR+D3XKrXVkUZrfVnjT4CFVoFXuroV//2XiKovO5WeeW1DIdeGF0+6
f/9arh8qKSjpRVp2q5VPyIFIf4NtA2DLxahsmPiYxlRKespX9Pq5SSAAiz2XPp/hntqWbYGInd4N
ju7tuzmb8Ci9e2IjgQ59v703RlGHbFjxLzFqNyvVjc88P6os1Mjm0BB2yrSpzxiDp8pdianaECJV
Kp9DQSZwAMm79qOlk+q4k9NxU9zjKAukoyNtLu1Q149m5Y9GhYaVMnhk9EiUmEPhOWEIBBJvcUyW
7Y5uR37S4vy7kvdro8otU6W8a4csKeQMF6syzXaEHISIz+/kw5OvChGgd0FZaHHTJieMKtJALsB6
NcpDacfCN9SH2zLTjDpBv3iJTOzy5ZpIeqqcHErWY76oqD5AcDqQx1YQ+vUk3w2/+40IXR+YrVN3
r+Fi3x8MkcQ+OFP56RsxFobIYHTmBiy6f2FpPZvTPcUTDk4YitpZoMNKBCDLqVyuskc0Pn7Z9HzV
mjwcoo3tFvWOYxAP/pJxHgrmr8ESe2okiSq/qHevlTrYy9CjbpXjYHHYh9W2lTLQ2zU2rvCL6+oy
Z01sceTAUmlwlh4xaHIvR5tWYjadVK7W4u/gHPAdgV5E1WPyBapXL1y7d44NOt9JtN9Lwe+LWKdD
hf1EQGlVhix6e9GKw7FsBe81jFpr+Ey/Tlsqg7UPrjN0dJYvC0rQ10iFNhxcsIqy3v4aod86hhKV
oZ23PIJtQlw/f56qgRfCRbrHuSENNbA5sJy2BVkgLqtXNna2SlQVjoFNINB5vflOP6ooZ3WVLgpP
TK3fLDNx5HzzVISIvW6U3dwFIwV5eHp5NMcOmD/+gUQPpJ8zODmtM8zQixNscl59Es9MTvy53Go+
g8AxADVBkxt1dMipomxGiXgpMdsTThkHxhzeI7Sfg21QLkCVTGuazUqnnK18NPJ/bBksMFTFNFXe
zosdQ1yF2ZK3dPIMwC7VZGDxR+XEzkDpn36imdGX52YD3t4ku2MVlJ6mNLCnMRgfp4Ls9Pj32MOw
SuGUMAt1gb1spN1P4mofyEW74S1Nwk64NCIUsZpcFfw0vF+rSwD09JO1rWkuiKGMGM9azchqCHAZ
XARzHpmG/7ZkLXSnJmePC1JXqd1ZLcUYRH2S1oWHpofW73vQnolVRgy7soTu8uTBpA2CMpDSX8yT
SIslMALp+Vc/xKDGTZPaGQWatAMZm/BMJnUMcZbAaeIrCzl/lgdC4Yn8Q3G6rlIrfeBi2ahE9T/A
BEd4cqeOeeUTOgscafMg8tFvkel2xU5mXkAQElL3xz93KtscI2vMkneoosu77kPgIPuju6hpi8vE
rTYcBq46j0j6UrA6Cq5/WxvK8WZFDZAptFVA52tA4hCl26MIngBAjafmO4pJ+/bzqmgVc8HMp5b2
RqzzgZUL/OOZvUJMtwXbPC62z14HMkDObLQuNRdM7gw23naHOZOpRUasFTL/zi+Oo1uNUioc39O5
59Sa45LSnaAax0zZU6fEa4OexMqlt2prtDDFvvQAjDUU17y5dmQcJxQ8+VsGKm5I4JpMnaqUm1AG
H6MZSt/BkN+pviH3QMCeePvwd0xaIoV3uQ6yelRBGLdSSo/2i5Sp5r3+disafOJigfU0UaVFWrGz
uORMTN+2XEeJeRMlo0TkKz5aZvuvTDdvEqhaOL88A+BpO1bHVqkL4I/OmWcmOgZCQEhCIl8KkueL
pdSeeu6rdBbl5QiPpG9Zm4vp46mUCpZD89Ky4+jkqe2kQoVm4OSrJl8kcX/Jc8mOMVT2OSSKzvYR
hkDCntNV1feEFebaAAElX4mV8jHfS0/Mgpg699yxdubO4XZwkdaJ4OGyleqkJFrKlY8rri6e4nLF
dsUlXSJu1+Kh/yknoaXX0+HfrUuYC+JY5fQksfQK01XdelqMyfvoZ3n1S88TAj/OBJ0wVid+QMuC
18OgA/8zQDUIU/nkiHJbQjzxCyUrXn4XL9uUfH7L8OXhyoH1ynB+qe3nwIj2UOdNgVwjVeWEg/CR
3fLlsH9H3vnHyBIoakBIMPdFlormEDOGECucHQ+g7ula4vCUskF7RtS40t4HT1J6lGrVrzHQKywT
f8wzlecE2J0KCPGfu/TCr+jLbcNieXpxA6dUyuJd/RRwrm8YK/DABwen27Q9hUGIXmRy6TAGwp55
/2SEJMBt+uXBAVriNf0tEfCX5IwN3VUWf93ENZ3Kuk7jjuLi3eIr/oYtDU4JxkyPClVheLQu1Caa
xdTHuGNzDFh6son1BxOAVBPbaRjv8agNGApLIEGYQ2EUTtwChWQpObb9nGf22eDzv+++TnKx4shb
HBV+Bj6z8QI3kb++Nl7O6PX+pdPhQiGrmN2chPAIfQxwJe2t3PuAL7KPslcPc7ja5950uwWoU/4a
Y751agDPhX/rebCKKaP3bz1l2YE8F3dgLoy0wI0Pw9LfAvaSaOOI77vDXWWJAAvdAd6vwKmqK771
HFLnlljj55nViqxD6oeyGANKLX4MnGiFTFJ6OwmsABIeosbayys/6Bl8DHgmUXkAzkBGMi6EPaar
1a6kM5gvFr7vapE1Yl00zL4XEViy3JbBNSAUobKhXmIcNfqTmlFtuA/mYuEPpgLUaC06iPpQUwai
mxppHMJ1inmJvsJJB4zn/T/m93ZsYF97AiXgoOUMc9f/VzF1ETqQWI1mxIL3ku11xZ7fH1hDk3us
uCngSxxEmvTdstylGUdCSmRZzSgCsrTvMLkHtH8VClr/xuhWQ5Zbftuli+BiBgMmCzVeqUUeAEyN
MzrdwkMHuEKdKyj4gFSYfdfy8UN+4CjIaZy601OSai2/2j8pZil0FASyzs/z9kR3XZ1k+XH3BbbX
lUJgCOROgABJDdDBkP4ZxJBw8ic6csf0w32SmNX9Jv2vX7del1Bj6Cn85yqxkil7LfKzoKGGe2IT
9eao/l6jWlOLbqMw4/DoT8xxUQzAc3WzkJhEwIM+8LTslq4SVuNhpgMrpCDTML8kxJSTLTa/5qvp
4jGfDCF3NkXCztkCLXN+v7Tv8q/BETE4F+bOZLCbJJ3nUTEy4TmXvnici8CrU7CIZc66HRzpuM6r
ThoZ7OV0gD24qWvLhdUcJqz4Qy2YSnS/FMv/3tS4Iuc1Aza9MlO9epMcNhTKUiZMwEiOKKHX99GV
8vYvGsUu7ZMgJmgazSbL5+MV5ZSQG95zl8iMJRgEY4iQGtChISRmWMjRPEibjN2KTlwxPRUX8UBB
+LL6IUPSIlp4eBirMzVNNPFV/V+BeharRfuSpY6tCaLRFZsJ86ES4dL/q2KV3Bz7YW0rMvPysvAo
iZ7HbGxFEqlQxKtxKdatbwCVNYf3yxXWzkUfdSM8jzUPfpz9oFYdJ+fNNX7A7bUo5xlb2hkAO4GT
Xz8ERKUUDK0U+GwQabGSqZ6txwTPSIW/xxQlJPfEXI2Y4KUIVvBR3fCpi2PzKgXBoKMxERbTxQur
rbuhVmr5KHQ6fps+yiY6iCyIieyUfVrH7oSaeeiYIF0QdNY+KVmFBzpGHz30Vj98Pzf0E3yoMJim
NzRgZUeR/F7xiVMc3ed0phW3yxrSfbh0/nKG4xfN08Rp6vDkSuC3xgKg4q1g8ST4BDhoK7c5Bhst
/QqFWbQW8tgerq7Q+qy6RO5z4h/h6YFFMLJSNodf87XgpBshSftXHtT3HLYLpLSyS5B7qhKpk8JU
WQbecSll4FdG9kx+pdp0j0hjvoowsZ3qJotjhYJPGqJCPblorQ8SQihrLjgnj9GHjpmKlOJfeX5I
ksZDPPV3POpfkD3dEo4KwOaDtchCbZqq7m4gyYwh9Bx/bSr/nLzF49WEG3y28YUNDQwEhRQ+iAnm
staScrEUpUeHnzpcfy+xu5ZM4DollBTimmuSRlOAbe/3Gh9/bdMkLiIatsLt7ZrBwBAVAWi+PZv4
D1INhEI4GHCXfffKGngXwnP9Mu9Kc8RJq7Qb1lLG1523qPNoV6hXeZlXvacKfw21s3UFGlLhhZrV
Y6w2ymugIPPnTtJxgGiGG9pV5yEhHxxVsmQ9lQUabACjnORnkO3A0vnhJoJ5g1MsrfEDMG2UBP52
KXBe8oPPWtmF9uSLIAdirYaB+mbbDXWgff9KE6/A6odsizUXS+pG5wAgAJTcyOl0aT2KDSJVGNEF
of+WrbFa21v5eIMQPEkV3Tbtzqx0ARQvwEsugxVM+e3k39LGO8Bg8HgQ/aNAKdttUeTUsoSw6Nqm
gGW2KAEPXagB3j6qSjtOdP8a8GBX7C2+we04efRIKwKNj+9SvPPs0solW3s699GmiA0L7f6iAtwy
LaZZm8hGr+laN3tjxCON0iZFktAFFVBfjuoG8PSr3Vc0KN2WHcj3Ka0QZ94dtHrjwdVaqt0dnRw+
3wY0C14tKULRgNdpUa3uvtwxBEAuBNkmrbe/JNwwHLxUJkenOuM3fv37E57nExbWYoFeFfYnCgFp
BCRtJJ/XtX7ZdRgSkSMQDF+F/hZwgkE/WDslTGeQN4xKGPd8Lc7ROJSMSE2b+ArOq/Enr1VRhK8V
jiuFxbYFv/i5oL6/5OSD9aov3rQYKilHtOYD04yxz/0SRT+8FXe3P5PG5EXr7DiTEl4G9w5TpJI9
5YCxJsitnBjYq10nDt5jX2GueOppz9KlS2JrPvb7RmHZmyeFJI1JWLgo/kYzq02mgjdZz785nRkn
54oWGF2jlnN17PNrrSQ8KCi1JaKiVo+NOD6LhEgU/CHcMvGCXt9biJZemyvRWiG2RVkLVAvBJe9L
NTWLhCN+ejbnrhTuMrJ4juyvBLcP0g8LXJSHWZngg5cwiOp1pkHrrgOWuZMf93pj/Q+VeQQa1Z6H
itdmW0GHidaYqsRzfKyd0koxLTPgNUoX3LIaioPWZqlqad7RaTQ+laetG0t1vdMf1VRfzQszTZsg
7F3Gk8YnO0QBBy7EES9p+7fnbURosR40Y0x4CXX3+IQXc04bXodFwlXgwYjR5BS9R/Xh+A8y9cFn
/YEip4V5NwqwBP4iS44jrSOIgbgOo43BFI9Wq0lGa26fBCEjBsGAePmEl7QX/Vm2B3wffLG7TKQX
94uzr1Lk/3b1qLEhgJcT8HTRehB61XV+X7KSuRlYt5rZxZqRlCOwL/WWBHw13jVh1rAlwkNyyDvi
jlEW7l6L5/j5PcQ167q0GhdREBf+XuEG7tUn2F1MW5kCxuRxFjiO0BGrdAK7R2aRogOEGxvtzR9z
qQ7QaLEe1NFaiVy/NW3UawTgmkJ9GB63zZO1nNgoiPDeyQJlJ/ytA0J8l5JTrmP64K+oZZKt/R0z
Fp4z3Qf3nAjK5GExT2mpC8oN2RnkDXU9mv4fd2iEgo07XPuj82G+tEogs9JkwI345fxlUw7SGGOg
aL3C7EJeQzWP04Jn2IPEH+LqaHN/vsiEGVFP4u521O0lFkCOjaE3tjnL2P1ZJoCBQ4MGtefiRobE
DbM24/Z77kOQuvxzvRyDRUGEktn7v/fQciInpLNo9ypdDtUDOuOtfUXaj2ro4VLsfX5LBcnnccb9
Bg8uSZxJ5z6g4ryKnce5WX04lJLynr8O+NWQfvuj5zHWQKe3mmAjrbdB+vqOerE2JTPs5HXZVHdh
TymW1VOi6tLPVZfqJeG3f+GNXMtvqXTa29QQuOjkB8PZ0qjoDUQbiAIQ8oUK9GYujEKS/dZKYR8Y
mKrV2iQ4PGYMkjyvZYx2/4pGJ2NHNczIBwYF0LI8ESdkMI//icOK0JEk0bYfAo8GBJ38ER5dPtdN
S2rqKcyLrvlRPvMt2jq5/hJ7vFr8ijjv16anLzxb8GqQMI/2RXXTzKcziW02rJBu1mTZRZ0mnWW/
tj/JJpJThqytVGu6Xbe9c2ZYPNi+YvYh7avFd6ZP3yjlxQRyr+0fwU82VCl3sFJtIP0joxNidupa
DM4HH3lOaEXsOZqN81l43HRXn90jDdlgX6IRMUnXLxODWaqCMal13XNjluBQFItPOhur6YNU7Elm
hBTtk0iglmAeqAUtCk2hKv7M5AVxlI9XTCbfFuXV20UwHPGq5lm3pDirogsxpfe4TdDHcxg077pV
b6pvA7h1Sjw41LOzkb4Gewt1UkHPjH5G2i7NSCj/8rOhN4EIHqjD9+HANuNmng34Q+pRdt1DPzHN
Ca1IVOxu0ezSOw4CPzv2Jz4EthNewZXTqnIIZ/N+nu4vNyJZQOvYXnMozWu9tLA9ZgQB1VaSf9q8
SW8XNgtq6GrAWR1zmluzP4fsx6Jl89YZTPZP4dLNcLXuGavipcVisrFSsbCLzEL90szizlQhzsLO
EMAOUD0CVQd31wDvRzpW07lak4xEJcQdlKA4+NWpg820rtbxmxInMyOaBUiUupS858pUVpsbxyWf
BgCJ9YDXro9gVUTh4ftl1TVkyaYyflHfinkyeZzn76xPOTCwOk8J9m05ugs6ppe3muKWAdaIDIPb
9zzS3HGAPB9ffAEPC4I5UH1wW6HrNHtuahAaw+0Pzg4Zu7t5ZkY813WRmquFq4rJOsCCEKLJ7wy8
OqtilCVkO9BBQbQariNb6SMF0XGw4B4gSYH+gs83OJTNnXtu8fAZybJUxsuQKQG9sjeNFAUeqsWf
pnW6Sa9CWuesKQ7mp621RiuXGSDUWFHyMGWDbx7qBufP/y2IgYR0R+zWgR2XIgke1+4hDkN/1vmh
ht+R3GuDHxr/G32PvX4ymG7ttywy+ImpEjTbBTxYsw8USJpqmGTrmeDXT6uaIl4B1KEiVciywWdP
Fex0Bx3876OU97ECUeGyoR3q4q1PHKcowfY0cyqfjZurShVsvIZwHavQ1vstL4jsAMc7lExXUb12
ymfUtbpO4XIRM1uRGXif7cgLsnI7h/8lXTlkw7BRrCG2irblu7Kme6f8u5E0KOEgjq6c2gB8bWW5
vTvRSUc9ludfZcMaNFHj/A65JKHrOtSGUzTi3lQkxO9bbW/8ZHdgS5ABQNZQqagqpDGRqUcyFXxF
p8UtjV54wNrRVJ2qx/b0Zd0XKRoGL3U9iURkTqDl1PlHRv1XZ1wijnvCvWo0UyT1sREmR/NlO+De
sgPmBH16cDG7MpXGaCdXFqsD6Qmn9jkOYdUAgwEwaIpIXfvKGbX+nplF9KImNai/yo5VQRGrxx/I
cyFW0eCpDWPTdq/2DSjMhMG+oS7hMAEs6y7qx9yzlU7csKDRTSJDfl9oMG3IFUHTw5MZ+VwhRpbd
j+7G68L3PlAhmZTKf2wz02dUgRM50BIwjMrjcEOWBfKsYkqy72wVkG2EpK3tCMh8uoL9tflc14Tt
TfbJ23zCciXg1Jx70Q3Q0AQsGeL6Okp1VwRzEgtepi9aFxrLScWttzMWQY1gvGpTmROO9GOrcDFB
DtTEkhY5dfeFwh66vm3ubzxE7kFZ+oapUjHlN4c9kZSzeVizUYK3YDVZxpVVe2Er3624txIG4qjo
SVQfm+WSFMyMAgq1Oedv5+6Kl2MBXing/H2gsaJmBhCsyog+zfjbLlWw61H8z1frW098sysQdyQ0
svp5YVZDpgho1tYRa8/Ixk8dk/koj1ODA3peTKUo2kx+0syOuR2I2oPTdzIkbuUhtJvg8x8Z5m1f
gOzLAQITE7z4lzGSKOF1T6hAaZtJJJlbQXy172Spc75/nKPEt5w68xDv68uvxxPbIkukuBlZFCfe
fPgnlZ2AObeRSEZ1dv/HhQgKrsYdCpWpMU0Az0iqGsDrd7cWMZxj02WofnYi2TTt8I7y4oHmEBTy
B6iBOh7eSrX6AgmG1wK4V1SFy4bhYb0u8sy0Y+z2TPe3596QIiz23TTjf9j0HWz+GkiS5O/kieOw
b3ip0D51esSIqGrbiLGZzuBb1hZwcKQHBEwOytjolN2lMFyw6HbptcCn5nVHmvw6TIPx0DSzyzdP
7qFo/hTpRlRWJXz2k5fyaXWL/4rW9lgzDaFuRpylj2ZgbZ49rOR4001gUdRpusHS2lkzHKVB6w39
GlEpSp127qNvnVYdnYHYFB1/bUmAnWKX+esMLdwIbTr2mrZK+4ldCC4Tx+YbpfsvEdPaPx+eevlt
cWQZWA6GXvEgNjdCZ3IcSS/30UBU7YUkeqyyHxi/pO3Sp7FBQ+CIus02ESPFmBbCrt8PR2pKFCLl
rwn7QuUH/k8Vvp75qGdYAo45SE+NlFrmKEYC1Y2kmXcs67r9xp2zsOu43L78AJ7sLJUVxResQsUr
0VfR/u5Jpgni1DU21oTpirAoQRtTYHv5TcWjobq/zY8WRladtLZvIM4FaPW+wNztGkfAIDA6tTz7
xpm5Id4U6ulCWz5eJwi5WuK5tt/r2JrrjJ6Uw4Ezxl+THJuyT42/zH1RHASYQcRycXbkOAYzzFA/
SV9elDKa0ocRXHTPn9H/gAt/NkfhCTGUPtNxST4VFL5lH3tpL6n2OQ4izFyr2+rMsApB02/+4hM0
+T1va1KUfF+ullY1f22m870uEOVmmcgl6GtM8WoihenaBMenkIK+Kan9RxwqjjfnvgtUE4OG3PZd
BolwEy4cuyt9hHA2fVIG558YV+tBu4xSggrz59ekwNOvb568djkUsNfVVdKVc1S7+maNLdG4gxsn
vP+C42YTghIgNilGLU1P/piDReYtuiUaYGqf+S57CcEL9hI/qpdPvyT+C0ZHyqpW8ACYrFOf1A91
E4RDPasLCYXXD9u5CMFEUbHzzIvrb3TpJlTThRgzg2XuFJ3rKthPQXDeq5mbhSGvHSAFC4GG60yl
0J5C3aHLjbSjOHoQuDdJJxZyJslIDyDuQB9Fjx3P0qofcq9HiswqNqzpCHiwFTxm94ASBU+DX15v
ReMiOEXxuj+xFKlm66+es62IILWopkuVz2Uu5zKq7yTMOpXTfRSEyHfXdjk5qokpe3PWSqxnuKPx
bSupQQUjBoOVRdRf+cDZtKfHIf1WURgLwkouAl2R9Qm++62A3tcHcxOf29YcbZ+dy1CbT1nbSpMS
GIIUtQp41ZPuB5eauALWUjPWvSE8XKDGwp8S0uDYnVsOT5P0FBTp6gg33TErhXJd2ylcXJOrHAW+
WjRYY9YsiKTnt7Jag4iISp8pwRrH+RzDlIUjAJemioimtYbV8LzYWL0LAAP96pMrH1jm60i4nwxk
IUCbK9AvFt7op5TUvFKSopEZKEaz11JPp6nbIko9I6xQGmj0xjWjJwKPTaN/XJKEtitlgIm+FWBH
5fErTDinWa3uuFLX4hGULk6y06I5CCpGoEz/Q512s1B1d/lIyXTTzoa9i1/T57sZJIdphindbCT3
pOQHJ0kkQm4/Mt+HeITAcztrJm2o+PSv6OAPlq5+S9vD0Hi4PmbUlfgcJ5Qww2vk7phsPRQlsle0
Mpk0xBKc5TzBFROMswbpJLV38DSWove/WMqb0A7cmW5GCO92dUXxTmqit5ImBUWgyeVHptzVtGUI
3s/z3KHSQXtLDqEkQwXUr/nlZeCyuIZle32bLxSgiJoHNPnhCYBrB+Ha7Kq99/MkFjTBvHn4OgUE
rFrW0nr24+BOWGypkXQ6iL5ohANXgu9D4f7rLMSQ8qb9YioCiFYjxO74i1vELufc6MraC2RMUV2L
X8786bXyuJ1g83vIUjxAWGJDJslMCrBXJdcsdDbCCYdUjfM/qe8kXiflxaHKBahXemtqe27Zvxoo
9kVKid5DZobdNldCglVyKpoEPtBqd+54LhUbmFijbxCEvC11htZhAAlxIxK1NLpnSs2AdxxAhf8D
sUyLxkSGr9nV4GhwltI9EuGmBdJ9fhQp/sOsfCFgawnoaZqTWMPTA2/8gY11zCkT9Yk0L60Koved
dD4bqlHBrpjIMVTx6VkVle30MNZu0YEBWqH8OEZ8g5pVvXwcH7xXPbWi38YOFnpfttRCNWjsIwth
lk6NYARPc0vI/FMJUHRCIS7dLDt0Qih6bX+3fTuCH3HsqdQOIIpQkzw+j5HgIY1Mec0jXXuiC+QT
0AQ7P/1NzBhPe/NBIhHbaiA6BbWIGvVEJdJacebV5VRU29lvXpb9ONBk3apjRNU9cCJjh5ZXE+KY
8Z6Dp4L/HJ6b9IcmzBYhG5WWOaDgt0DDbFm70usu3i/zASMHv+4W4ivcciIMJLXtDaOePKKGnZBP
iYcw0xZsQ1NWhijkV5r4tymPY3FIUDAuHV60QEMSLWTE2nqCJU2ovFH5DWRNC42juMe5TgC4v8zu
x8k+XknVv+4zZ/QWHyA8xqLJQh6hVNJpiSw6HMC7z70MezrZLLkO3xsIHVtuff1qsww7biQwTCMH
B9UNoruzpt/18dLuj+MlatsB6Hp3NFZxo9owUIdvumDsBuAJ96cCDlsBVE8tc464KSN1D1N99pQr
BzT3Y9aCxMt7Kkb1i6234iURddJ0JCMR2R3ye//I0Lpx4mENhMKDBb5Fn4xbhuA/tHn3pR+ssxai
ZfFHj61skIXVpEU5y2Bvw5Uo2suOa6tzQs0YN/B5G8RDHds+YF3QsW8cdffKkVJz3G9GgGCWWN8m
Q9N/ooA2hni4ziBGOgLMglPy+bFOuqnnHRpv6k8faKTDICOBf9ja1GX0xEUevlQ9coiavkDTBrwL
+a6jn3YSEY/iSEh2NNK/ejPTM6aP54ewkoH5wASuKnQpCRnBRRvezZEtpALvHje62x6QdeTqEipS
lQLvU6MqrfpNGp6zYuNsxt9jVNke7mjxjlHApmMMiJ2RdyROLQ9tc1QrrOQ0VWBy1J8Kdivi4tk4
6inlbeTLCbJ9SubgVRYIM66Th0eM/l8r/sIau2WHYWTQj7DEV7ia2r1I7fKHaCqfOYZ++NIS71Hw
kiTUR/8bEbniWLNMQqAdwE61yYUhkIk8lwtSd7umgWSSprxcN+m8SDpQQj4ok5/mpsGdhQskpjZ5
T9iTvLBjvQYeBaqP/l+78JTRsLcMtYjOB2DHtG/fh9iyLgK/lPALnUFS596Df7KsRNja7goAkCAN
1o/RKDXLVDaVoZABby1YOlZYgTDDEB9pbLgWOrk4V+HAvL1y3btzMILAaNJpO7QWBu2aMhNa1zGv
Bl8o3MMZ9Qcc4t7+0V8FUKSGwPOZJKg8iUObVEYaRFDbgc+P2XDav04f9UEk7X9uKx2Rgqgmeg5Z
rTlqF4hFOZ0aaatiBzRwzweOYFL8sfTAVtWHzrObhp9+yOdiHSrY6Qth4CxXnQgdHauBNm+nnYQA
me/PNMCs8OGg9/v6LO8Uyd3dN5oLpAnlPzLbNgqE50KhoM3RsvMG5eH8cUjQSKJm8tWaTz9eJ1Qz
U33h0VTtsjsZBVLPOUxDJe2Exnp2Ctu7toMtdH1JEg4eRmcl7MG7ul/qknzuF4YT3XxZuY1BxOvu
nmC4zXmJgYeQzoXPqf5/krkhZ1MWWaU8m8Mq/E/C1oB880eauDmIH1DZVMIZqNlHBOXEYNCEhNfC
KIWTMs+NZRwvXdlKBlXnuoFhDRVoiHdTN7Cx6K2pN3Q3lQwWxJYWhS7E3APo+S0vK2RYcUhxLYrC
wixmhxmYed2E/O8zKQvSTxbq6hI9+Xp/AtJtGGFOdIxG/2RjytnC5BvGc5Opw2Lvu4D7YlwuQtab
ijedsnL1fRduQpjziLLUdIO0ENya2bmap/I8TQf71oUYlJXFORUOOj0TILbLrb1o665QwLZ3Ioeo
Sd8jcFsXBaXTZwmnBGq8896mpqjIpZxSa2jBN4gHJMNuGVLZxVGCEjQ7PjOKTKj/KxlppDzmJdon
veWqB/ooZNgED6A50BBUgi7Zorl82dR74WvKcS6Pu/S92Kh8Et3zjO/+MgAcpFwNUUOtcNI1S2Zr
7bZQohpijW9Ixxw6XalgjWCcE6iBMJwu2IK+E1iDR5CJ4IBJ1TTgS+VKKasDyWImBZoJyGyoZEEY
jcCTRUXDE6FquneTIh7FPhBL2Rc4sLzrXg6KrR/oK09LFMS2ENWX+ObngAMiKMHtvyPGltQ/sj7J
u9JqVyXZgK9Dw594KV8TRnGTTB3wxmTsDon79uMXJHznQFpuGqWFTXU9koJ5ilwoTUZozvDOlsrC
JS1uxSi53Axigkfp+mq7YO8Lz1fZYmZ8/GZNBYVGT+v8ZSTgyVwc73MCi/zfPaXAclewusucfc4j
YmU3d9OdsYEWzRMqGpq822z2t2Lrmnk/iwBYzysjL0tZ/QFlctY3xOMtA8Wv96ew54N8EnGnsLRj
EC2TH9/OAxSj07eRnhoa40zBhviDt3keNhw0NwZEMBrpH57/d3bdJV1ekIgEeJlVO28g8YsNZMw1
tm70V8QnFuTrkg8r0YQ6Gv24eic9oFhbgid55lINdrM3VFZIRdnO0G427FZGMQmcMyP64IpnoxDb
TTGu5uXjOerXCgJwfSZRvJeICY7x5FXXLgVzwy/+YF16sN6gTV8kf7wcbE1fzVRZ+aH3YWcwFT7/
5K9WxvCTZuepSNp9IuszvP4igIwgN6UfMCSvH9XioWuo7/JfFjajGOHgCu3RbLNSuvzRpQTXL+N7
iKBK64vR9I75xYKrEg71yqxGwIvdpU2RxnxDhKxs3fsCLPkonCyM2kX/4ELKUdYAc73srDVB7aKZ
g7gqpuR37Gk0dWlZLOSQLTdZGULG9ZdWF0YFFdK2QE3BtuPwWyrCpVme+aEnV3sQJYTSAquVwu6U
TAhakCfS1hJn4Q2oNZXn+WqdmSgh1JT0oIy3e+aq2cDoTT+IqA+4p/Swsbla94m9CxMkAp5w2oN0
2IvQhYDoAMal8mC/wPCeqgjO6zmtI8KOFtck25V8Ok7e4uSL8zWOMLB9ijpVsWORk7665LxX0BHJ
uRXhVkFY9nL4pmezRZ8lqbS72K4SMevuZr63bM8si59R/HYKaTHapjZOr/QYU8EI1KbdLDBplZAZ
t3yToqnrAZqiOaql4V3C673SBYZb9v3Zmbpwtrf4qJq+CKcz7dlrFy6WO3MXmACAo5g29RFd4e4V
K+5f70MqIrzSWjkPUkMZ/QvHSDI1oNK1T8/E6B6rEok4489MejhYw1dKJk++lDoBaJKI8fAxgLdU
yIHXlp9DcE0xJY3vIAeYpIr2nVZLVht6VC7mS56+sWvgvTnmItrkyQzVDfIk1/owT1ThuMFpnpCo
h/Tzk0YrQYY07gfF/IM+WNm043NcEe2QpYNQ5Wa93s2PJhk4+x+sb3s7xGj2Cp6n/vAL2ui9NQUG
Sl0PNgJcjM23eGGXpF0wAF53UDVJZW4gDd08jJ+zR2bjQlUVEHUk3E5uS1iistzaUR+x3jdNH4bF
5R3shlteDadP9HvqqkJRLGodti7mefnhL0g5ALePMfkr1bd3FJokHL8qXcUdWAuQtmxThD55N+Mv
wzTnlZBnRAZKi0fDEA39ezSxikM2crw/FcuNtEaXA5m0+Amskrsp4KlZV7Awg1zcy8VVo8GIhnw/
fsVWfY3L4uXUMWIqwfvxG0Fo7eOifW/gtpiRwNMcdjy9oqwNGokopRGnOjwSFy68oa8f90ssNQw7
5NkpaaY+jhM4M9iqh2XObJYZpOHYOwcoD9t1k/1S3htaX7Ssi3iNM4AYdtl5KgiUbMvIAmYtU/iP
/3UpbsjuSFGSNQ7uvFcigVm1a+EfaYdm/m+Q/P0EYw1t1Y9ZcPFNlCbZscPKuk5R5wd9bh7J8FvI
li4YGjQuqfHtxPWxVIpQRvOtWLlbuHnktEE+L/2dryD0pfqdJZt31WbGSYc4E1F4mnELknI5ZQc3
OSHG2fuFvb8sOoQ4+b8egb8GwuGYo9+U8VOi6hxViwj9RSTNdQdPXhzqQZqkoUMVVuRIgCoVSU5f
P3lhwr4yB2nxldk2uRZkBuqZ0nh+FQKVq0teZBHW4U/SuGzVpxvinABKr2OiF1bf7cND0d3oUv31
WgpRHMGuyU2lLqnpZmAHTDZ6JEJ66eEcqzw4yuqQXA+yXS0X+HRWi+/WWkjWrhE9lEzr90Epd/Rj
sFCpl635LeIC5/dK3weIZG6raLng6fQfnOVE5QyZRu0Szx5/25oyf3Z/ru9yQ+V1y02W51f4vEcD
geGLxhpIPF45u/XRfg7G0kQ/Bs5/i666DKt3ky2vaLFkoZWMeQ/hs7zaUlUjrNFaKv1BHnEXHUMP
jqh8mf44S96zFgNLbJDb0zFsEjBkP1Za895LBzc2TSzO+rZUO0Z2/0yPr/LvTWAw/aya/kUvIpVB
uOBzq3/tP07BwRIwvGx3OHIlZGc4VOwo1H7YenhS8glwO9QT231YSZ9CbEgrgnfQqD7scgoFqLsv
PTS1uG5wPgGYlGr2YyMZ77lI6DLBh1o25YlvyRfW+ahBWX8SfC9Fu1p8Qmh3BxJgI2vHBdNV0R1S
RM1JX0s5nK9B3lYNGvifk5wBTxbowgPBbvBe64ZbDpC/0f4g3IpX/EZUvg6HLIw+w+ULpe04D05G
KIkO8j1MJ6XzW6QkDbRhvFvCn9DCRMPKz/109fy58HmHBEalPQqRc1/X1gDCBoDgdh9iF5kOSKZZ
My7MPubyQatIsELxaoRpgf0719pgqtvYXSU8bFNHkpCAZHxFESeXvAaGn/bEF4cWzp3UBZwSpi7D
Zt2SwXfv1DVfjXFe6ynO7gYoivKhhEcIImYzWmdQCOXEPqQjOyD1/WXU1w4anpXasdZOOnh74Sau
i5Z7jBb9N7vLfldH9FOReuYLVcaAoGfyWX/hii86ewRrm8yi/YT+4Pd/jvigCA1tPrKIblrmcjXC
CGaUevQTZ6oFKjiqi8tZfslL8vQ+wpNgAmReAeYtF2/rrnn9a/qzrgP9/tJ6BBS6fS7/yIWYUnOQ
YZ27p7xsDhroRLs/JtIIm/fR1ibFgRkmXtbF8hehYvQ0zHFNEYgwq41cMDRMkw2jf292EynnWTL7
D9kI4+bS5uTofK4f7Dv89fApBVI+iD0Bjrf2HnP2C9QmD+OpoXhBqTBvunxqQIbHszdfHVvDmG4p
hMg26VOwxva0MCPh7OybJ3+Ny2G4mgykGFUc/SBIlGwVtu402yJEO3xdhbvKF3mjuJdDa81vo4Oz
TDqe6lxkIPUMPDvpC1/ODz74IjnSk4pUM1Z7HSJ3A1nQiGoxnhLxz8/079PG+mP9OD/EvD+9gIFy
dv7pr4HEtCaFK6ycVgCQwOB2q5y8SglLP3dNLTRKp9KiU1LXapxITf/lUyzfR1KTW5E3Bw1KcSmS
BfLawpFiXDJk+SWGULjoh6xPGwBsKZ7zJeUJ1iXxUm2pdK+xWEcnNvzeNJmWRGNqo4/AhDP/W+mI
xGgt+FdNveUMzPQWUsDwpWtXRwh5MLJjyr13cAx3nDiKFPYVyd+Y/kKwD5ZBufIx5jI0uw0gATGT
7uIWxC7XmbR+Bwf8BF0pe9Nlv9aa7Hd/sQxrWldr6AFZ0hNJXkyTiV3YImT3lwg9+OM9wZ7sJPS2
ek2F1ErpgkP486+FYX1Kfyv0iAnpjwjs7CWptr7JIrw/EU5DHlC4v/e+T/8r1BituDclnjsSjiZC
adwTrIJSsbQXKRF5LvsvpVG6IImLQaHeGpfkFNuxVRV6+y9xdYlh9xLhG/jLCnCt7jJH+pepiNV3
6UfsIxV1mE8LDaK748lsHZzQKaiMJU7YZ9xjG82nytu2NWBtouYZqyF+tZcq9CLrToTi5jDs9t+9
rVL6hZSULKVczaG4KV8FkJJrhlaXzI5/EAidM5g13ylmHLwf2o6A/x/53TUniO6PbXrF4MTEp+AU
lyjbk9kHIsLwrXsGvgBtRPp878mNae8XTdfmrwDuRpa5Etj/vN/A7KtVqVEVwN+5TQQoGGuMC+di
HJe7hCGiALN96SvhiybhefnVYJEqrrfSKADyEPQSv+HswP5wMBAbP89HoywbrcZrKVP1br0s00OI
/65JRCKiqkc9CSCL6r5dcQE6Hn2JtrsZh2o0IZZ9rRa3qzzUnLpCYhY5OjxHBuwOJDaDD9Qwo/W5
dO6KSDCi4qs7eo1n9aU44DmkkcBR80lEuPdN3gxoqbTPbOazBM7Hn6MtQe4oo3sWKME7iNc/mV3V
5WaTxMhv0IDpFNZsNSF8oppwB26GyVss3EWtIy86ZSgcfJOqDBqEEmQw/YNGTq8lrCkCSDILvh3n
k+MtmAUKcPDLcniivJvi4JtJHQIePMS05HMorfv+cSWXpAdcXYhxuF37z18oVQj28Tx8tzecsm1c
/2PgphSbRDEQXx4+d9XTivSHWDVmpPkpo4cUIsvfoeCh+7KLYo3qRait9Vc39HlFBfWVYtccX89G
jMMvDM8/hiA8N1cs14o9djbzze4bW6KExBVVo6AO26dSVgyHIFRg0FoKOTX+Eze49ZGnJUUiaBzE
YWYuCONqJA4rbEL+XzK4uDqjxozy4IkH1Us93rrHxrb/r9F3zkohb45k4hS9bctZfkQoDgDYLr/4
xV+MEUj6a/VuIYh2oQ4HwpcLDDCOTOvpUBwWWo8K8Z20heorUdwy8Z3ir+cwWSqiw+dK6QX4Ft6x
CGJAoa2s4j6gCOhUaHUyMxryE5FhEf5Umt1Q5h9owvqDDSRLAnw8r2g5SR/d8wfaSSNzfqn3flRp
sWQoRO15vByrYj4NWI72RycVQNxThdzuOTxjk7gF9x55+ecZS+HPAX3nfHwd2Hlo9fcBuF6DSZL3
HFSBWQe6hvbsceDyvVOhf8E+ps3ka68cy6hv3PW2k2fFMgBNEx46ypxeqt9Mr5bQCk31cLhR0S3V
ANpGccV1GQvytQcN/fLZdzePJexdyu42XSLflT7MdGrIpu+A1ukd1TG42UGj3Ihlxu5tTw866LVD
n3JZBksK17WJ9GkJfPWOwdIFCGJK0jmDVYT3NPVzVbna04x3qnaarNIt7KFPp5OKJdEuPEH/gMNb
LaT3G2PzfJtuAN/YPDC7TBLNp8QoraWyH+H/JYNzNI7Mh9Z9d4UrEFa2kQlh7ybiRY5Hs7AmPRlN
wrjVUFGAF63lhI3tvfSX0b8mlJ+IyC70qa4/eqYtEPbdYYUqZZi6MjgxcGjOWxRv0uGiitu5gIko
X81iQi8XcCK3y8an3sJXjcz+73PBRvGc8jCHxLmpgJGmUyyYMnSM/Scym00TmCss+MPIW7A24k15
uFY2lGVO9VXdGnMPOmuKOMqH445wUeEg8f9xdAl8Xk/5BWqkLN3gsKhMGyjgjAJp3JwXvAuA/ScA
FBNZ6BLGo0eiFvBSlBj9SJmueNMQwuv7DxUP0ag5BcI0IDchTC85mptTWxz+mgN4mhL76URKAud3
s8dZ42mVrtAkB3VR9uNF8UuME2IDwUuocsd6Qki+eosSatdi784ELrH/vdDelMGZB5P4hZb36hGK
5pOORXH4O74zSvX3HOYtSjG4r7AnsDetmCnITjHtEcPln/bja3Gg5tAl2UYQMdeGXDrPkexxTbVV
BWvDjiAZtZKsh+SWe4+TpWOVNBnrLctyITCo8FGrEyknGcagefc8GgW7+1rgdagVANZSwjgh0pWr
uceSuAvaNunKhwocXdDI5bG0fAtHmMT0YUkcewO21BLZ24AHIODeDxChbT8e/eyDDPx1MfL7wGP9
xJhmfZwSHD4wGsgmqd0sJHlEsVgVi39cArOPKz/uNmhQchsWlBeGGpePTQAoLKhXQ2LgxbUtFkof
XhGbYdxlNdC6fGLhmQGwzZV6hQIWCvWs7VDQAPJJA9NZ5KpxhGEEwY4MBBp6JiBpAlkfKw+8Esi+
ZoS8S15Y0cztJBsZYbw1g9gJeYwDi9ygVt2GZ7gsnpDzXBhJ8S5+Tsm9P2ikb7HdgpInkCPNUs3o
UkpnzZSlAPnejaGzCmnIpBkP1TINf1hV3wK4M8gcozU0imSL5/MLjgnMtcAUDJEq79kvlsvHbbF8
IG78oMDrvOV/rtLv8uhBCFQ8Lxz1wbGduYZt67vGYPhSSc1wNxWPYiDrZKsmbH3ILoMPQBKC+Uu0
BV9S2ZzrKYtgjoO0H5IpwcAH6aypAzYAm5cSKzEw+IBRr7OvQT7Mc6c8WL5IW1AJBmUAn4NS4IK4
TcQWn8Zk23YQ5frog5U0MgyzgdlLrosVTS9WBmriiE5WiOjMvy2zy/2FABd/qCMWoILE235Et/tY
7MF1/a9LUYq7joYr6L3uSDq0hfUso9mFgPYFOb7HKnwBSnQxpB0ifNEkozcWMzIzSxTRniyQTERH
hecOp1D0n6nDFfLmTm3mWCeHqShkxZPW2rSTj1zVBSWgdqk0l8qG7aAqpmgnRfbn/6BDzGtRcgVm
DCvieNTdp+H77wUq1Ed+0cHNZa7kF8uDFRgPD4LWMmKepclD6DfaYQXDi8RhYvUM428qrgp44Gsd
zIBrz1Ci4ZwOY+KF/rq6I5Rav5V4AOE2JQ/pgd65kmHeqllEo4wNg7JWSK27G1Gv6nsVPjHxxsbt
gUmOVn2bapqCSM7QRL2huMYTbWvBWs8jY3uzivgaeF9xt/+RsgCeBDASlTKOwkXHEhSwi0E0L19A
B1gazcYZRkfgziWM4+khD5Q45drwBWr5l8utKYUITtxOCNQByuvHVgbuGAMDwls3yHXDF0xygLzZ
7fdxZJpoVLcjHhXjrOgKFeonBEwqpzTASlqUJFYwuX0MAx+6AppmcEQlE19UIjq4GjfgRbLwUpwq
2Mth/i4MJLCu/vaSsrcJdhsK+YdL9xH/yrR1QeixGLUwgiQxHffWpkbfMTfh0EuBaIe5ihR6mooj
9nC74C4x3jGDpFvokxGvyh8PcuVa5xB38fWuoWK2JlXaik1TOcz73ZCdpP07I3n6I7EmuAI8eUx7
A5QPRCDRIDon3dBAFcl++KR8Zia83YbFUMQHDGc/z4l7TjTCLi1BnIzW1ImnIN4Yt49mMsDcd7Pf
HdjwYA5szR3pBV8NMzRoNH0ClvnHwotB1nSTQ3v40JoPAv2/KefwiRJ6QUPStoDU7Kup/8ljs7NX
lozgJs3lZ+ogkBgWn4EKdxrZ8Efmqrj8ERlsYbRCxqWTrk89E4UJP2uIwN5vSdFMENJC1lw4SIxb
X82DMh5e6zN1Dgma8YdD0WVr7NTMiMrkfqX3nT/V68bn4eCDQNOiDARB22tuyRaTyUJIhMrYxZc1
MFs6FIi/v3OS4EqkvbPWOQL3zdCFAzqclALSSyPcUY39IiZ/wxz807mMRt/2IPKNiVpn9HJXET2q
sU9WagG/5Zn2KY3cMc7v8FOhc1GuBadLLtpiESI7l9GZzlEja2UdIUuWbGA696slhNXH6f4iPuDH
aoUXGUWeGzyChETesXG0vEqoETcixKglug40dM9Pn+/jnqj5Mg1+3BJOjK1wlDNn8oXH9UrDW30l
5kRMi5M0ERqlCCoIoLKnPANG4ANTEObTPtwTJ6AvdwnEdu1xj4JejnpVBp+CXy/Q9LxTbRDpNyLp
7eanigvJFca3TI+udsQVNq0DqRLyyx/s93grhBxclx4VqBR2aAGGf5Ctp5d8hkT1iFgqNsos5mWp
MylgRY1viFB4YTDtMRwjrep1J0ieRJHbrjvB3/w7DSI+xLENyCF29+VOX7cMMVhlj+yGu2AqtHRY
9APLbUdJ9OKRPk+3XaVvnqZL9/u8zl4xioxPdeKIYx8QyKr5HkHl7eGUATKF08ry2kHPlR+KV+As
ypnf8hNTlE25/dwEEiEwC1YDy5LTUPJymobvE+DDrHL9si+w7kADI9/Ss/+utIr8Vf+yZZ07cNbA
IJ30XztasH40iLjXXTp16+5BC732xWizKVLQh0Sgz8P51Fl1GfqL7prU96w6gDLIlMFwzG1WWwOa
27mx6ii0xynksBUy8ocwh0E/K/04ehJN+V6S3mipPodeyLUCXk7AMImhiPSflIJBntRKIH7jXTqO
d12vSkRE5SqExOyM4FsXYCAwrcgz7Y11KIPd5Toj/mL8vHvsOJjAgiv1zb9bn8KY2oFusEjgj97s
Y1w7x8AhJgQ2BhS71okg+Y6vT+jgCjtibNek80bU0EptcGx5paWKmdQSr317zU6PDiJnfGzikDai
73pS8KbsDMrEaNGvTKxY7cTjOPZG5gdF8sv+u7J4qun7xUQ8WwrYc89TBfbCrTOQ6S99DUB4/cG2
BFQd/T68M1eqbO+6VT7O3OhRneLpylo0/xeTtePgnrU8fiAJY8RvZ63U50qk/FGeBhSmhJsmQW1a
8viMLybXeeBT7X/T8FjMPjY5rrBVLmFvgvPcj7WTj7XIpPmj2d+zN8jtTydxV3NeqRV4aBt04uYK
VpB4r00WUX4ZzcGKd84EIjyOJxVdV6v9SNxYkOq3YJnzFjfTqfFPtVYlSTIxL19SABrAWGzmHj7K
d52j2EdutvZeaPntSjf52NfJhvhHdw6z6dZrKxEUtysyVqkpZRKIcXGPb9cIynutswJXyzy7Dcnv
JsYsGc/zjIP6jVpwkViUc4BNfHLQHij+AAqKSsl+bemDqAf1PiBpA+5Rzhy6mjydZUkfSzjfadzr
jQ/yF2jLRd84VzKOMu8TLBoY4kW62MvS8SeYavVpivNDj9Raf/kTi28sNXpJ6zD1iF2IQMn1vNvy
2h1PQkUUBsY44zX3iwrY/5qlyTURApbiTnhyvBvyCGoEAdF8p/xoCWt+FU2K624iwXhIQ0fo2pDF
wfC6IIzixCu1OJqkp9ZocN6FQ0UqVPFXEvre1ZRNwjQLEigGd4mHSPhsFjzMBPLxrHc3y2BtR24p
Unmdb5BlJv/sYeCZ+PCpaLmi52NpP0QOLvQhFbBlB53OSv5B+ubHSGh/O6aS6f+U9Wu9Qdm5SnUc
sabBuFMxdHHb1bFU1UfwhIU2u/oZX0J0yYzgBQRQSWLxWrUxTpWkWvUzUuojg30kPFORszSfn80l
A9c3Zxx3dUpWb2HpzxXgl3IjC1coojckSeRFpMrUXvqL1Kq/isZXPLx5F7QX1Oe7bZG93R/Hecpy
bVPw3bvYr0g/ZR1+38VDnfq3XduH6F/VETUV/+6m6gf8lSIWtl12QzniB7oV2jKaSBob6SKva6GE
mpNsmaRR2PQbJvItQijsWd/Ja+Ib1kBMScRIxVlexRkSDFVMC8WB4a6BYs9a+JmsrvXtBj+3YWsy
5Y9aZ44N6QorBXzyejvmUlDdME2ufhZSY+022nw7uA/AAeLCvt7ukSmndrAC90W3uygCxAHtyJml
yLBH8A11CvcDCUobXe15NSEJLIpq0ZOIZhOcRa72oDkar8Lz5gAWE+N4xmyR72MkED6KOWdzDM1a
Goz8gdPRPeCqNNJDaNgiN4VDEItx5r+rG+JcpoMZsMQuQNcv2r6RkajuUGotXShnhmBDiR3VIgIo
LWHow190u5mYdiZbQJPAJpjZG8ju1g/FMQ1XFHNEICAfjYDg+6+g/NiEJA0dFLnn23kETmtVLlFn
efseMU82lyBa9X6c0Q7W2vI6XiHWr16icw/ku8kPn7zgbiTAu2kQpwtHPEc5TcwyQpZRQ1c6Aqfb
HjBt3MQ/jWqFBMLCowATFRcLvFz6pxX5cICKOua4j0zJDrvHrMSNM7JV6c3L1opwTXgfCE0K/GEX
sP05UGkDUAYqhstg9hMlQccyRQGkNgc3PNhEWZhk01l0t2I/2VeAQ22j+DjMcekLdAPyTFXqe2MB
ToGqxBUFgm7FKio+Ac/qL+qKs4B+biyC/75sENpOqzZ4hOmc/cGEOwtn+i4D8/C+WigSDyP/MjSX
oznYKAjRZg1a+4AQZ4kh0EuURw5LzKpnH4Upf3k1irYzWpqK+Cbl+4Pq0j9KfDwA88audAYpdW+i
Jvq8c9DwOPaWV4Uf7NQblCjvi2mb/yguBVlkKQq2uMHHSw2Couz0ztD6RPoHbT0uq/nKaf18oGhw
XaNPqtLRkk7W8Wk+ZVv/fNKEStClsUannN5f3Kyl/McuQFi7o30nf25mfLwIFUQX3vH1TbRXNSSE
YKMGOPINQn1sQGrhDFBjvsrGXAWVSxC0mXtZrXOS/fsEEl8EezBt+miKkcfBKRbgHAB42E6iF0z2
pL01w32lDoE+VJEm7f8pNJP/S+7ox22HFrK8G0xdSfaGp+6DM92tTc7V/mllL5O8aN7a/TOvcRH0
rv49PLWvkta1kniXUWaKUGfHoByIiUd2mLfA7ZqC8qxR1YnJeBblX7TlfZmKXH3xI9IT3Q4CNnQ6
48ZewjAp5+9rcgJdnCZ8Lp2ZQh+2fAaJFwJyPm171ZU/yduJUIrl6WMpLrfIQmMFUY/yo+dOiKH+
Fv/tPuBZz9ijJ2nvmbT9Dfans+fSewB5cLm8ENvFMlt495I+AzjT0MOD6BXUMfzoigD3RQ/M07/m
e0h7JZKQX5jgWeOcmi9AK0i2Yj/ysk/OjsMV+w++IS5lYWPd434filnHyDaRvHGM14hrzy07Yc91
NLNr+EWbYid49THwVOnka36R1pshVV8Xxgk2sf592LEkmqdc6sGbf//PwKjTRImsJJsCXu888wKZ
cb257whcVb4S6Mh0XyF/mzd5dL4eEp6EL4Mn8/evaoHtpoFu837RvkyNL2pKrpCfnfLHU2fbCi34
mtJB7tTF3FCIohKGVWh8BF3DVL6DwRbf5VqQFmASNc5+DVEEXouk/0RwMixuoXA4ieVunvkFIQSr
55vFm4cUcyREVtwMNCrfD9/cHVxDc6PaoWst+S47iMEuf7KlLgU3dGX55twYlTNf5Iqfbx/wSA8W
wTdhxpd5xYrcQ2nq/USqEhdHna9llnxND7cZh/zn32tx7ZOhhpdq0hzentKsBqBYrZmqAV5UTATX
gZTEHqUyO4Vccl5e+SXDCGEFxHKDCIEgnTC3zuk8nskZ/+4dYgqh7YicGss7b9wyHtPH9CszAYc6
FtjLuB6xA8FVQim05sP5xqxqNgkrm7SHLoNuGhAFUJtsxz966R8fWV6DN30kPSaUmWKNphzmYLOq
D/8GMDLOH12SvUd5ww5OtBzdzpDln4ZFy/4B42wVOWfL0qwqS3+8LYL67kQ8wsLz02WJs1w6Oryo
8PZ1Se5xcFxGBds7keugr3m7HSaOtIBdNm0u/53cRiFjOyBziYJr5eQQVLjuL5wHQ16QyuECKxJG
SgsmMr0tIl1hIKAIbnI8sm2ehVRHHHXKaBhzIrgwDfo6b7TZlgyEdRer/fZ5s/3Z53Zot5QaKTsi
xKQcqNkjaLb/4s6brEb6zEJ9uh+AE79j2Fl3uyjCjWAPtImfb5F5kzDPXzyd6IAlzUtM3oLCWoLv
WrGY8IYxv7J9pESFP3ykujmbpMNcdXJd91N8EJORSBpep+T5+RgSQ4h4GmI+ifZIj4ET+wUoXg+N
UqkGRNL91kbpjiHp2G6MmMCeMnHnfV28Q55lZ/15lP7AqeSVrjJM1lDZQClBwDwjhOmwMtPbxrqK
Ao1QIKgR68Ipa991UMeYLcvx7q47BDluWmCqii3W/nCFhETzFY1AnpnUn+Lx1wcmHk9BBNLUisOk
RONjKKgX5YkRw18mMKodFMV+YDlONXZ02Z47vSHAxGRQVI5Md02b5/m0D/dPXdnWPHh8IvC5HK4D
w3imHnL7e87QOQUhmUaW0avR5O323bPeI7Gu1+rkTdUwCLWTxZoROphsH2c9WfVFPtYGsEybcmaN
t1aP2NO7MtMd+jVgnvlTY0kD2qyzxllqbqrXO2E2uSxCsumCudzmaBPtZKkIEQ5SSuFUOjc4uemt
SjVmv07mCBDWI+5GiCgfccEerjWboaH3ggVZWBXYy/TWQrV6ogfTwRdV+0Ji+SgeclWh864SXM/l
krW1Z5ZrDi7oSHR7YHN8YmbRyWJl1dJCZ905aaXOPeQOtFjwxTmxFQcFABTP1iUoPYxB3LE6MARK
7JwjUmbqvs1mW+adZkj59nD46xf5koZFIMP1Kk5VDelbZhpBFW4L
`protect end_protected
