--
--Written by GowinSynthesis
--Product Version "V1.9.8.11 Education"
--Thu Sep 21 20:47:36 2023

--Source file index table:
--file0 "\/home/cod3r/Data/Gowin/IDE/ipcore/DDR3/data/ddr3_1_2/ddr3_1_2code.v"
--file1 "\/home/cod3r/Data/Gowin/IDE/ipcore/DDR3/data/ddr3_1_2/DDR3_TOP.v"
`protect begin_protected
`protect version="2.2"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.2"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2022-10",key_method="rsa"
`protect key_block
Y6h8cLpzueQd5MOZvCcJ5gxIgsS3T4mutV9kQK9qyFnV843dNquNOHCLmCefsgnWKEpta/7vfFL/
nfYQaFDnIyTao/EzYARq4hjRS8n5+Q/qAJV1CdINi/6XW/KHBTzU+Tx3V7UQumEDZYTdWcamvkZR
w3siM1p2f9ybhkLOJ8CL+IqU2XKB0Z02f4M/1idTQvSZwTYQzodGzA2uPCauG1WmYwZqU4bnRuFg
SoYxjckJx6ESLbOxOlQFLp12H6kHOLq2V/9WKreZ17m+d3pLpZRPsrVhbAKNT+fbq7tlzBkt+4n+
HnJJcyV1RjYwko3UQSEdX4nz0OXWtTdY1mMh+w==

`protect encoding=(enctype="base64", line_length=76, bytes=599984)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
MYlhClIZNhBnFLurri/3T/Fr7qno9AksMVWXhXOigs8P9nT1afdw7nzUVcOALIKw/5/JuywCyeEU
yI9I08sP/Qx9qjWIY1HpEsdtRvxMZ9gUlP5jatOYdfk11ztcHxddeElPCoMJYDqKItXqiOgBt7aa
lyFpVsGypGg7ZctlGYnIYS7g7Dk7wPLCMAM7B9y+a62y5FM5ZR50PMfmAdd8sziyVpka08yjIwxE
PWafHojYn+wySrOl0MYj8Jvf5hJvv/87ackvLA/nHZWz8GYGDdwZy2otxrNZkCxdysvA+AEEaupZ
zWhrk31TNjsRZYM7BIJeWE1pL1o4wgEQSwjdw/duB6GlxtYyUuUT5EkldVvVAtM5hSq2iKMwXegE
1VetrhYkWuDEfVzxoare4XtrB+S75FG9xL21Xai8qUcOJc8GvugT8+LNNq0wsZ3J+T8XVbxVfzre
NjyqMGSbbj+wLvk3IQpd7kzDQc9Vxe7Ow3yqBAPUxOqwKjEpP6cqrPrCN0a23y9PL5AON9mkOOKF
XT7J1jmS2d2MjVXoyrpX4XPb1EmL3aasHKKthmjDNN2ddwcMRA3hvx6XtkD57zUz8zolC5k/iQP4
lkGM5hGXQR2CvDjpOVsuAQTNHy5MZvooxKqQ0trpx7TDd5P/YFctcvVgzl1KjX/kkW2loOGveUHo
b2Z1WfTqMFX34r0IPde+8i8teS4fqLdB3ZQQ10Zu41XcBQiwwtWVR2pgUtcBy9Q9LYf2qCAf7vau
FwBJIlgA4bqo7vKdzRiqscmxSEQXNX/2ut8LsSnL3Rzu2ZfWbELeCwU3PEdo+8s27p6f77YpgG0h
U0evkrZixeE6j1QQpHboyaw7hJfcjJTa878hSePce7hl1+lyfaSO5+CoXjMF7NC9+jXoIbrKaaHe
yhbLYy4iVQBzj1sL+k9BbyakD4ROrXmFn6K0gnlOZitNFDej8vqRmL+cz4Y6iHffZmUkxM4w97sb
WIGrdsxvlu7LWREq2p7nLPaWZZhPR95TrazSd3PkI1pYxBa2y4xr/1lkUTWuItvtGerDUb3RdQQS
04DhqtnDyA9SeDVKYsR64U6Q8vfXraFJjJUkYwSISsEKr/Zk+IXFzV6A/X8QfC1EhNoCZ3ORhz5r
XKADFLMsNDMAuNmSPXHdHE642c2sEnKUuKEgLLzqouWidy+WigLkL/HM4xHJ6a1sBDdNvnTEHU90
FbK0QaGn+9N5dGT19VXyOPzhwxC8X4KmJ0GqouEKAufNapf5EKNeWQL6sC74IsXW+bTD8SxqZLbl
gA3Ao6eKpbORcV5acfIUY2jfqkxURGmaiHIxeY7RgpeZMvqYCo1yoDvJ3mgHGjFolHeKorPU18xz
iwKgi79ef21WwVbp6q2UUHS6Rx1YvjWRNBm8B1xyOz1+gy7OyX6idxNwUViDSCKgCP1e3RJzGZP0
xN3RoOJ5oQmmY087DlKVMHbc8tErGvqOWNwI1dLKLljEst9+DXAH4kFJBPVontmynGXX2WTva7s+
TjY2pX0rlMx7j1hIt+xZXEyG3GUSIvoCOFbJaKn9ubV5+c8rS1kIvjhvX2tDKBogsXvKOL2onh2Z
lR37cTGZEBygVOOW+9GKt1kzT42/4Ion1cQN8rpZy22wG7MtKIlONJveCgMxOeOrjqeriweqCug+
HgENgPZrFHGXNmMbIYgTGRrUQj8H3myJq26zAhx//1Y6RoQKwDl2aWdmkMV2mXOk/tzVQsLibTyC
9cOTv4a6YUNJuucEKC+04sjCfEkFBlfSXkbMgpKntvcWCRGY23ghU5w4IFwuiIILwfdItDR6QMNL
3uE84QLFsuSL+Iynd5EZu3gSAJvyTQSL8miYTOqYRUMqQ3t9779ffqXAOOsTRcWfHMPwwk3M32hr
zlQnPmuNRpmtaZFTeO2KfVWci8fLPwWt0La3dYzAnQscArQHCfNwjgkJeLGZXPezwRN2q7Wpfzbt
wJbpW45omY1MudNf1mbmDU/G9gz7AWUmZ8wHJJIKJHF/cjqqOL3StT6ML0sjrzg370ScbBPYD+L0
E+GJp+CTfhBphyNTXQOZqG6droJ2Yk2jmFpfJHk9Cb9oOxI2vLgb4U1cvtgsa5QnT8c69tYAjL6R
oAbtehBd8UQxeW7mdSF3pX7omqlUmQ41EZoPLaENU3EC940OrahBFQU3JbTXZUJ2yqTN/bMOlQdc
vH/BUE7yZQSjuNYpqvUtRLz+SAYutiVCA4ZbC3aixLBvvAd3P7Ke0ACiSESx+D356QFUcir93uyT
bVf7DbG/eUw5UbyGNSfnfFAfRxxAZPuo9rys6cep0zlouTL7XanxSYbPaN/NRZsCaGKEsrW5qnnk
QzZrB3HsA+lA0AWdlHqnT76Yi9F01jUOPM1HNGvc/72OHu8B75shBjkunubUrsIA1gjfk9k4/Ghq
D2JjADS6F2TbNNma/k+RtyKTHasLaVrrEguSOIkZH+9MIdKhvOMUJ1/d8oLhkuIQZyQL6yZToLE+
YfbgQUYxiETrVpQvZG2DFEfSpinpXGOqdxys8e6ZcaX1UmJAt/p1Mys24zOHgMNJSPMIp+kV4a1K
aOGAitzSH6jfpYnyjv9WneJ6pyT5e2V7XnEsfM/MZJIr0kjMKsGeS0kpWpLVCY2niAvMEop9hz6d
D3AH3/KeILEL4UFucW6bl5uamDKL4GUgQIBDALR4oNH5PerZ731ZVCk4hFh2+LU+cbXFuH96WuYf
6RNQLBQ7/Tuc+XjBWVry28+3ve0jPbohusYWk853c7baWVd3YqR1J6MTqpyYILkUVDrWVRX8gDo9
rKuDjs+hmLm+AyfZAz6T5hDDMG6CYB5fYN3kRo4qaWmROQS66RLromgMvjsaFP/kKjYnl3Ggg5B3
SlISgW1zrSd/jJ72Yo3vC37K0qjO9sbEGbq6ElZG436NWbEdN25Busj8L/c9jmfsBMe+0veTpy5b
F6lexQybz0Mg2MlmkkNpm4YzpJ5zaGfZZlaw041Fsyc1VJzAqHKjSb29/An1/mSEB2HjaT9dWeFG
8rfdLdtRTjnPLsbprbXIqKObpiM919nl4Aakcattbz0KMZVmaGh1moh0qYbF8i6fm/hWphHqaBrr
7LjBlRQCoYM5yE4zm4FC+UxAHgongf11wc1Oj/Wjvqt9+qCjQAkM1bHhJ7dyjpCoJ5rCqsbwkSjs
EhQ0ibcd6K0NeSZRBZc3bLr1LXA06Py7PFWzy5F9Iy0I9Y6jpsvXpMwxkQncSW7VQjnev08TyMTN
YhdrHSA3ahLOhTcLTMgtjIYqcbPZKqUeubUaWyP5OYbTlCKMIkj/45MIo5VVEnIoXYlEZ7Yzct13
94nuneobtkfIN2/IRNtuQZFnU1bmIf6vi+NBMifNXbq0uWY8y58a/fc0PIp4QaJ8m7hharzhbic+
o+HB1HRsZMRYysmZShi03H+Rg1awtVRLEjgBgUgGEaD0LbRG/lqKAtkEbmL9hK7vT5NhJ+t5o9SO
ot5WHB3Qukd7ZgYm0y6/0Ai2lbmovhM4F6LRvjt5HK6dS0uhyllLB6MHpi9yPIJKkh0O8Z4qgY3n
6MufpawWWBglL9MocVP4sULT+jgRGU3qlKlbbQbgNFwLrLkK8fktKNXnuvu0Xv4e7dWFKdX+6g/0
TGjhPSQVSboR2dv2EzzjuurnuqJ1dfkZcdvJ1k5CK/BIwTQbDZ+QTzV76lC7TIj3VXwSNgABQ7Ee
eIj6MRoFaUjw82Gcl1nEsXztbjFNDPVUiqp6PetdoP5t9JIBni1CIfjKDr/s0O8+970UPmrjeyFV
0GCHx4Ej85aLfgJDLKdN498HXIA6KUj42HxRQovSpY6qh69OgdszKHcAzf+2LYl+8V7NfXvAkKeQ
FD1kx62C7cXgdHQsOWIsIOEbyTULmeUHUXs2f0ZZ2s2TPEkJWhCoK/jiUjV8krAs/FV4k875GnA5
A09s1GFTjeuprLUBHy3v64FFNRR+77SZbFeiL6jMSx3RYpmh7tJYM7Ll75Nfp8dCT0ny3TudzrhH
S6UBp1SnVQt8ucsFS3nk3aYTqVrkK/EfTbFwIqLkXZyNhlhe2FSXtkYNPRSd/rFpnsqA3bn9WErf
KZqbuLbt/piM5E7G01pXH9WlykwsTq5TE5yRaU0fBaHjCKBQlGvbDTo8R6yWC/XA0ZKleXdaR8zy
q4jsSv4qGEUh/LR+TWQs8AnhyeJ/geVwfHqhcGQ87mVVwedqXgKoYMnaPXpaYoA0sl96prcvOcqA
645oRnpu2PZ2rNNCcAHGB6HIPQPK64OTnwuPP+1sxnpY9AT2UiegORRXADRlWS03zJwcrfS/USpX
L+/gm4uPbV6ibDJpJrDmsjjQa5KUmBI5VkqoNP+JLxpvThS0OdqfK9WdiN9c+VIayOb+IouC3iSM
WK28PJjsTc2t190qLACEwxUdDHRfGqvf3vd2Wwx/m9O/SCJS07k2hBgWf4vOKWiJHdAG9OlFtAr6
gnBKpNFsBfDulnBSXZkWd7+H5J2IidfwFxdspHbQiU8OmB6Nv7G+wA389amfEBJRF0J1dZSM0NAg
api7g28lcdnN6Ht+QNook9PlEfDEJJjGbLKX4jq1Y6PM88R4rz07DWBNTFz9JrNQyU7nVx2VQ/DE
AQD7S7GV0GUM1/SGp0tgbrtMMXXDb1L7BR2ZoHDurpgzITSvW0i4Bjz8tczkY5xZs9CWa7UoR+NB
yYaEIKNy/VCm+nlxPE8CqCwQFozg00d5kb2tic6bLwqcWLa7d2e1LfgMmSwQVDB6rpmUQuLdT7zz
8gWCj+tyxcPmCSuAvWUS9nDCGJ/tQjmQcN/BkT+sxwKKdpqUK1/wUcZgSYfzdsjVrVbPlN0CjL9c
4tKubIcwiHnBoVevFxUjr+cvETswElmNy7WNDnLS7sUBWcTB3b77uj28e3k5qhzhCJLNedmpxtnK
X3DaiikgY/rZMJ+ohqP4QRl/RaxHXwAehYOxbBYIDGfGVLjiaPSIdLQIvNWekwfvHrObafKaIUNL
PjTjfqeUvKR7KAOvRRlERQYgM4KCPkmi+0uHvdZMJ1nfyeFZQOiupw+gKzs4NRpnwvoDHALU7sag
3oqk2A5phfddEpJm3DYlrTy8jsN2cp5PES3nCEeJZDF4kQtJV8oFG4FRZBN8V3ctb3xDKcnSVUld
9wolnxnKu2TK62hyNhVyv8CPDegse/hHEL8xkhHqAUPucNFECw4xjqrJ4QEHPi3yom0/C+UTfdGM
/29UePp6tSs0Mb6g02JjodN9NILfY7IBUfJ/tt4hIv47/klLb8t8wxgEQx3uuqCFICL8/JJehElS
Fqq0QaCKnG7G46x51wTGz6T/I6i8k5BgjKJRSwcy1i0XBUjbDDu9iEt6j9iaZffpuzfRFvCdQxbO
yFUa4j1g+tdhhANazBbhRghQmgd4EJYO9Z6S48AOQ/63wIboOYznJk/4udRR+jxOzCqt7e+zVysk
IXXqO2dVc7VbYfK8L5kQcirTXOgi5eWiW6Nu42nNNx/6QQvuG5I6Hwu4BcIjGClQKYiyg7nGAjSu
dka4aK5Av64FoQ7nWWQsDa11eVn/tiMXIKspXssvvkeBXsdDwKDd0GscbtayeIyR+MgFmjciqlIe
nCnciic86lA0KKVr25uNMILA+ikT9YvAA40EGDRKZPVzZvIuZk4zt9Ch7wMI9ctCMOASBSQndBAt
jmCCKdKUYxNVsdkZwTHkcBHFxwvV93409sixbUxIlitLAhiSj2Sh6GcB0/SnMhSKet5OKYpycX4U
Tpt0ExWGfMt/JAEmIJVLV6/IBQUknqlYfCRjqfnALmBwLlPTMhNp1qDExEndKT08tfI/HfJcdMNy
fQKvSNvRchlcnjcXHYI60mnzOZGMGUvNzAECscwqz+jLxTs1hiEP5sF/MZEAP29Y6g4OzM6ZKBF3
z49ltAMZdmsy0tqSHYZVY0MQS99aIY28j3d6FuXH4IkTq9jGPiNGTkxwqpDEW0FBj/uSdJgFezyj
ijQI3L6Ttj30eubV22cOXCsXjkpQfugiYbSgTSZ3sw/wlca95rWOFr+s1Uo6G9xEF2cCB/y8tf+u
eTL1bAVnjDmFtVidiB0V3KCal/SwhMS64HNNavRYyuzVHPh0bXb/RFTTZnicpZGwNG5AYTlDiETi
JYpu5DAWQY2TPjIVlzuthcPKxg3gP7TvF0mrkhaLDBaOURM7LRK9jyZpEIoHHUPjiZkGl9CpESL9
ERNtq10RNS+0URrv/mJbLzM34CqADqKN6TrdgDQ55G2wu9reMxb47DXDVXQt5a6eHJlZrFboW3jY
mvraCuq/icn1guu4r6ifTOojbNtmvhA5VsKDMtoJLhPEZutk/+LLCulBT0697daPZHGY+CF/RZz4
P2O3g3fK331JPxQ/o31t1CJSnDDm4Dg+GCpxa0Vd0GSsj/b9vsHkfjPbafRPSJj3bQXeE02nCEcC
QZSclI5e/eoFKX0QYdmErCD4isl/prhzDJJNUsv3tHHurr6ymjeGJ2ncqy6uJFDftdpx0lpny8MF
3/CqgGWyaY9x41cQ37AIaE1gtwbsuIIY1EflQpOX88gg1gGX2Gw9tuNfyGJf9AWmOslvkbB8yrw4
xCKJBcxIPwfcrzYwSq4xztRtHZY6zH6CQdX6Z2Z66L2ssg8u07oVhbBQgDXv+T2hNfGwF7te9zWk
yfkePWCIlh+ZGYdKvYwFeniFC+mcBGSXNC5GZcCLiIKXB3xUDcW2CRo2GNXb2MLkA1EPxgDAVuKJ
xenWvTzBFISagiHhtgX0bE+FDI8zYTAAEhwFUNMnfraxaGkVzM3Rn5Lg+rsbRs9pUdgfIJuM0G/F
4S0Y26ky+bi/YcJ+bUMeTy7/pVmuHQV8ml8LuWJINalWhxNGpJ0GzERZ4ucSVvzgMuLAJ94lxggF
qyBKrEnG/fuF2jhUCGe7X2656Uj+FSSwOvsORU9sBPcbcxMFLvFILb8vs3dltYzUhSFDiRAgoGNb
xN6G5K13+h8I1MY6FU83z5Q64wAurMlOt7/w2bR6mQW9c2Y275yLW5w5y8tXVYAOuPfpTudfbpe2
OWGo4s0fT1pHSx8xYh/CWmuFDk6LZsWPqywR+yLs7y/JrFniYT+/yea2/hor0C7/6jbdAGNAe59d
/VMHM0zIqLTj6TXddgzYsdC06aHrS1xPeMxFTyxQBOAykXhVem+m85iUmq0C1VjHUiOmhP2GkKXZ
TPayzZRfAxu+kqOFs/W7eQkBZ/9Pj/NBSlBUT3UGCUPhT7dQBUUj2L+Fa9jYfj5ZbWWfDRex4uRD
ILuC5fttJO8cMG3dRPsHuljlxWyk/U77ohXuNZmWPekv3hpFdnD8mfOd+jny8OoO+Db3uFxIcBY0
DUi+tuMermMH72s2TEaR68qc3pEt71ZXWqhAXRtXg6i+pH3XGDTY4wTJuhKCeWscX+9V99b6Ruwd
QLArTXXA3nhh0Yzi94H3J+Ka2CbUjoHKvxAeDV+7ln3LB5qG970/c+kj0CsUnkfGUzee5W4GeUHb
36rj2V3WDCLme9urHvbQ3Enk0ijuvPfyskMgDS6H7m53xLH/QtVuLfFWYCQeql9iBikamhnKRrqC
KHdj8mV0MU5tyE32X6navxDc5mQA1idXVLcbr3PpY4eJPD1i6fOkCm+vfOv5a6raayUs163jeW4k
kOyIbc+Z/d73PKhHJ+xz1BD2C6qZHbsiT6qyHZQ91AnkwgEafAxtQvro+4MJ4ZDKYTyVfjQDAmi9
2Nv/WpPvFMhQGddQjp1mU/52sLBoTESN27c/eEVmZqDSSCwJX6X9cIgqHoltgHWT2/WOzJj/AHah
ebFCzjc/rDslbeQnX89h4PN11mabEDXu04HqQE/6/dDnvPJR/r1z3UcbT58TJjOPASPyW8FLVkDT
mAyiBpRPNqgrfMjVZm9bbqSZs4pCm0vPoeaNwf0zgcgA85K9yXpyABUBbVhADuR/ZMn6FYVNecS4
wj7gMi/BcERVahxn3vBnPXB7aCyd1FnF+iJQnE+yYfffY0tIp9VakeT10l7EkxNuTBuy/nQJNVUo
K4JIhBDbOgnDX2zeYk8lAmtcWrwzUYidN9gi5XIk/1PPDVRw3UTmjwfiqLoVIBv0BH3M94+yr+d7
qBvrSh4dib959BrTTQZYYUiTvP3M3WhNSeiite2EVDoSuUuJx+ShVMgLEopU7a6wvRWXGSsC4hTK
dlEpHpY8SLwFVl/Btun2aSgs1UfxAcGuigvYjJXibZkZf/znV9TrpP0DKd7OEfX6+gk79f2UM8pd
wSkqxR3rMQmlR4yXhowNRxvvxrUmtAMlXzBc6Gs1lgUt1t64J+VjYZsWEeu7/PnXanlm2/Tuq0nu
JOGAImeFmOo8l8H/N2OGlk6sAfYVlTrX+uUJe6PzWkjdChF8o+EoQMyk/xlzDWyCGo/t9uGVofIu
IZN0SlG4/Llp2qfQiR06hB2Er5GD8GLUOmuKk2FjcRDpMFljNkQ9cLoROQd59PS2Amje/LQYYVpX
goeC6fh0XFyfTVoCSeACNYc4vhhQHrmZzennCPBOH0xgtcoIzu2hA7QvxBWOZhhlZYWzCt6KeNwl
j3Et/YxQKYnXueIxoHKPZsP8COYQC+UIzrDCuf5bDVe4sxQZUCaWixXndDBlT4EnR41HrTZyhYkV
qANBZoG0DugH2LENKRyEnmPfbSQxq8fEn5lSdhuP+gxFUXUvnxwvlbVxosIPTiKrIPag7l6Y6ZoV
tsEHegEkcHFCc5ojngK9kZh1BMSC/q9md0BlOKycQ7iaYwKF5uFJEh71WzYhscYWeQS9Z/4CzW3Z
dvTzlhQ8jmEBMTzX3Vb3bvWyOKuo9rajxiOZAZU7uN8INePfH1HOiAzUHiFTEu4Ou/hc17YJelDI
G0vjbJP06ISbVM6xLs22DnEm/dLmwTXDNb8tL9mDlbiBshBoZG4ZtN6mpo0p9z2AZ8Ax9z+H5rL9
SS1AwC/HCHWa+l/4FwtC6pOYUz6b10aWqmgHO4FrPDzw+HR3R41r23QjfXo2qLcnmPVMyJztSDQe
66AL04y0SLE17Xb/X/JVFVC/H35hWr5HLYaSxJ6zcWOy4P7QT3UkkHR2uP3QFhaDxxmr+GU5UdIt
4zhw7dXj2ii+hFudgAtyd4cGVU+lofQNMo6vurV5ysU5xW+bwgIXhn6CwrSNVwi7yaRcPqvNZXcg
zeiFycd/oMbtJm8H7KnGKxhz7DZfbOGAIgOusiM4kU2/RtgHoULNXwZPGrbdX/IT3MANss8Gr/Zt
FweJjjWo/3ijD6M16C2O5oXblTSTw8oTGYtOn8QdSV+Ci/94DC4K+X9RY2RGppNNOJhMOoHnBTCJ
w8W7g1GK/FR1GXVwUcCSTse+xy/lAbsCHPku3m/D49tySAxh+oTE6fNy83XrkFszQeq6nxLRqk9k
fo9EIvQeUXH9E/Mlfxm7LY6OuKDp6mN2cIs0L+CFEZqQVN0BN3Tz/YpfF3RG5z6rPPPWNCp2kc4X
OBJdmZeZATHYLRrll5aZIw28Py36biUfw9AkP4DBtPAt6RfjZaiISuyG8nfCpZfz7GyP34tTM8YK
GW9kE2eSVuD36VRDCb+X9heGS1dqcxLyi50k8q8QooCPhNkAjgaLAMuXb93Y4taM0Qc+mdtFGlQ/
YSftEL9KRvzDXlBeWfMX0xQ0AL4wl+vU09rZ+4+Y4qtB5/jkfB2ezzJn5U12+F2U6kmOa2UaU4jI
dB5apNAYOpRtjpH/EYBDqBJ05tLu5bzOf9dTsxfW4wTd6jk3eVFKxJHuGWQz2Uu4W4lb9gpKOOMn
I8RWPPmoQD+ZohrSJqwEogaCUUv2I1Nk/S/C6e0Mrxd/8Lk4lHUsZI56cwsHxY/oippJnAz7gQ74
mlEh1b7sKl6loYEkIlx5QkNk1EZ8nKtc3ZVA1BaMHGRkK9YG6jjqjcECwAkBQ7/f+YlqcfzvkTOz
l9Uwug/Yuo+J4UVcqzgfESJywK/VQe2ZrBiLtFe1R7EOquxgyEL05CCu0oIouCxYPh6HLwjjyxM7
lOStvkb8W60Vfhvlnsx2TGCofwLeD48k4wjWMyZZMQaRBaID5KHMAFzLkf8QuX61YuIRiULKjJCH
0d7+jRjAiKW8bo3+qrVKS+8PqlWCS7c/SRaqx98xzQ6o92Fa+lWRToi71FlGTaJTFzwg18shozPv
i6FaEwqjru2CeuE7OosxWLFdsMgjdERyc8SsCgBlSjrTA36y2h+g2xvQnHBC+3c8q4eEip8yWdLu
M0HYorFdEU39VuSkufZBwp41ej2wNw9acjJXz4Z4HgyqgfV2eCax6DpbEqiAvuRpb4yTW5Z2UTMh
Iy9e1Bg+E6/NeKXC+fjHF2MLbcs4FWi8G2VZazCkD2fPbFC23vUfL2mVlWTYLevcvdFkUIMqkjdX
cl9lZroLO1BJ8h6wVkAAByT1ZAkxAh8w0bCkBMgFFM6WDpgRvUvQmEHpEuYwuAqXwcLfJZO2qrBo
UTOWRcK+rHcCw5mILaBMTWwUf8dWZXoOWfoH78SUFGucOdI6m6CMu+I1kZjP/iqzhrN7O9NtmYb5
nvwAgkXQ9+imPm1J7fNI4UEU992QeOAQf4lyRRi6pEQ/gedVeDktmY82VjlLMYpTlSTthj3+dGAF
k3rKyMxN+/cTEQPkZrYnLizSysmR3RZG5dkTOO4GNu6tiSrZvN59FAzNHYsIo6STww0kGeJdrsQd
9HOQkNccRbOnryMVuHtLv3RpY3XQ+JyBT2thgAoUfIWCNo5R1+R0IBM3paH0JZgq+R/8sW/9zvV/
CKVszbK7eujreaR1UVyAAOfbVwphbsNPeCrIsxekNjhis4aeCbktiYOO8zErstWaS1ZE0X6jOnk+
0KXfYwJ4x/Q21J5tZZX1pFe+hRbi3w89PND8MVYcjvI+GPt/RicNQe92MBUjBelaR01E9RPS07hg
26Ue0y8GEx8/bUkWknu2OKEBoLuAxpq3edq0q5m6xWozSMEgWStjvj68XogFn3DT18qpFYr3EU8R
b3I5g5hkadPfxNAYoRGyvNn5sR0NUVR/v3HZeuOTig8ZWsLUdipEA9LWBQ+iBTy9QBNEvZphffN/
912zvjMtQ3qrdd4cbv42CNqBLqWTL2j89VvlI/pAN8PYnUK1lHu2/I16tEIRba8Ic2gm0Dls6Mv7
t6J6foJqqcMo2cgAR4t9ANGxA7NVF27FaKyriuQfq6gdWaQlfnk8+Stibx7IB0D4+vTaCxQwlC4T
2fUdofykwYV3FXOxxM2KRsODbgDxEceEF+6uZS067t1oOvpfkDx5Znel7Eb+RnM2EDTcO8xz+Pfn
FuS9KpsiU53wf74yfxjN+DNICd7iCNdKZ3cyHgREhLB3dIytPY6pOkjugcInuZXdmbCYKQBwRqZw
UmHUjb2GcfpUzggPlBTExAxdVntqNf/x/f6XPQGKloUn1gHpnd5z+YYTdpZguHg5WIo9j+QW3ZuG
n3J0+UxSfukH623lLCnw77rBFlhn6L9aDsuTLGfjWRnEGdfAcieUMrWPiwHhcVfN3ZpEh4pDvNEK
YaeSWuKVhPGBmAptZ1BWnCmq/N3EBkSf/UGFpktLg+dXuuMeecRviGjePOPBefK0s6/uiUgFp14T
10WrnuYt6xeS+RAhK5Z4z23TKzRNNNJwWnsbTwyLfEe0B15EcDFKwoEpcfeSac8DHbyZOVc5Ozbc
fjt+0HEvzztNy4QjMWSZ5H9qSYLC55knrDrRDYh8aFaVIt36ohvMebK0ZOG5f3dUyhGsATbwwLNT
pj43kgvIKFCked2SYsuR+oQZojLLd1ZokQL9qVyy7d3xA4HMhvo6TGDM0DLzVLKHeF5yskZGGvh8
7rNhED7nY9SxHPCiEGPJcRRkdST3PigkeqPrVOOEVqOawkO8c7td5sUuDunoIY/0ytSIkV4If7PL
lotCO1nmPn3jpOvogb4vjiaBwC8OsYFs4X+olvdubGwTu/J550TANDgmEokAQVhpsy86WwFt5Plw
LlBr+8wiET8cCveAdBX2za993a9vDad7IZeluA9te1pPziiZ1lEdFJ2qXsxrQ6n2ou6q6B3fMOY8
61BJcGMHyA1SJxvpFEJ4LyAchUVDEOvpMAyxcgjqqZyGjTsh0spaZ99+bC4otgBHsp+c5QIlt/rO
rdN57tIleyb++PZfzTZUiA19hguVq57yOVClm2YfZuWs7whUxm/62/n3MHclFgX/OGNFGMXMDM7I
OcL9Ut70TQcisj8fZbGNARJ3i/p5NP6iRRaHmoaz7ruimMy3V1vrTA8xVnuMwTZWgRkEKJr9GgfM
WlPcOR6ADW6E9vAmoV+sk4Ow018Q4IxSQI+KHH0mX45pwFHtvCR3IfSLDy5Jaebzw6Y+c8sKGDXe
lpSyGyT5034L9t14z+OljjaqzCziN0FY9ZnFja/cZwMkEf2d2CQNnSYxzfiRLtCC4ViFwoFwoPC+
l2sxfR+PT1GazbD2M5/R1rS4Vego4wV3gMUVGu5CbS0qnSk4+a2+ygFwO7f/KGj2kfPHrhNBcy3D
cKQGYkquAkFnbB7DFDYELNrFI2IDzfnoW6XMROQ1bVerJL/fwVCQUXVMbAcXnp2cvpIFfDOrR4Vg
svBo3Oc4OFDDiaOPolO+nAWj50S9vAvWZbSOmgatZ8+VtRgGvNwGjEIQ1xfe3Db+Hxy9kOzXO1RG
257idWMnQ2qcSJIBIaL5N12xM120QmvkZmp99l11mcGK4rWtBsaXj7HSCOxMRwz+3dgQBqDOmbiF
TJIREGARg3NRevh6aetmPcIJczl9uZbt7QPi3wjTDDsIdyQvRMhecBCAyELdltkR0I1GfNtt9+1k
d7gKlvqNQUFWUCcguNYS8p9rfyVJw9/KdOZl3l0vJ2+31K4N8bEanqcsQqFj97xpuqwueKUazqXk
vukleEfnYfqf8+IYA0Hyk5DNyz51jxOPB34FR4EHL1Qunp6QkkFl76qiE5zXPZjaAiACKXKc3KsW
AkAEvALtxefH/rzwNs0s3w0Wwe6bjcMoMU0/ykSqTtjjde9IjBUZvDwCYVbSjnv17+vdvRyIEFk4
gu6RifBDYiCqUhCWj979VTPHcdmzUDDXBj1acVSl3dja6PNjPwiXF40PRf7SBrtP9IG9rSkOk/3L
g8WxlJHHkwq+QREJ1eHg8OiWHfU4uViqnX3ncWfvAHU0CK6mP2/omTJ+hyM2fPT+PpCS7TQ/baST
Cg918Jss7btkiRDoODjCnFY63Nm0YI9T9lgO/i1UqNXhykpDyVe04PRZP28UGqwwFgRncCX8W//p
PHlA+ug2oMgodPRU1J9I54tGj+rQNy+gqWP9MB5mvHEAs0XVUDhWWV7Lt+ie5isHe4P+ns1NemvD
HdHE5u4LuTMe9JKIGaMqHC+YmMR1CQ5aofBPDcXr7hRIjDF+YhlYHzRu1p7qsS8E/ZBZOdfn1BCw
xwSbzEDw/GozsIJPAvo3PfZFDC9HWkFd9A3A2dLhfmwV4MU3QJKGi7sfQbFOLKvMfj6Oe7p2dRnp
+ziOHCWqzT8vDalZL1E120zlazpxC1zgKFE6vP/70Ph1sEanX5+SWuJSjaDBw7InDMT0waDwFy/e
c9Q1iy1yuiiEf5jEouFrl4cS3PPJnqNMX7wSZI9hFzIqdhLjMyx0VQTm8BPObGnfAzweSnqXNKkC
0QqXPw6rSYGTZV242rXD4D6rS6nBGzqflXI1va1iRoxxRShFHyXOevqBUWkB0VQZtMtQMLvIB7e4
uGRzlHB3DL8ZyUh1uLtY4f6BZsfmEqPQRjfmmLvWgDq2SZbnGMM+V+xDlXvfJgwLwhw7yKnMEk/x
4TXl8PL6n2Za3pwCj6DKyIMgwZzjDFrjs4EYmTWl15Trzzq+4fxVvCiRsg/k2aWHsW8qdRN7d9P/
OVUjcQTRGoWR5pUGaEDaY8ThXpdGp75emKqcQYH65iKoNTbtTCjbBm4SjSFFmX5qFJNIUJIY3MyH
iHysIJOC2rpKqDMpreA9kfOMijhk1MFM6x2CbUoBl1C/HXPnnHsiqKlozm4DhtjhxzqPWCFmsKik
GEAin43V3pUCBZC6cnc19jwJ8m6BTw0R42xkarkBHrNDdyQvMkZJ8qTngHM2EU++sqIiyQZJoecq
jjyXL2JL148IaUtMuLqsQ3/Nnud4/G46mNYBWLTJlbn1kgkikOkbbqBfWzS6ymDETHr1VgjFZxZi
a6m+mlcvfaHmK0bnpRqb9Da4x8ruLbYXNLPMuCTb03i3BgwvANSj1atYqMgXCOy11ibGFxZ+Cb1Z
h2atJoY1iWy73zqlLHqQCVa8i/1CzR/xbh6lVp2xfCZC3uyVvIbOb/37eDZljrSE6PQMIOmScfJj
cjy3w6+9NiJzoYCwkxXyo1HHhN3PAQFMvvgPUU4jWW4zHVvn/j89NNQmNTLk2ZA02fQO7icSF/SN
VrJrg8l8vpwWO86C7bKUnJJ9F3W6Xc0bhIaNoVRPFuR1epdqpbGZnd9WpN4Qa1/DCE/9zYd62fAm
yzn65NqwsiYU+AbbP6OnvPQUJ0toLTK8c0evr5SNEKYVpod+6IlgvLsx0uZ0F9oS36lqcRxxflI7
MmkrwtysGScl89yxmK1YS0wtfgRfHvCPjCkvX3LsnRZAlLI5gY3lbnJOub+W78p6suaUN/383HZt
+AMi/GGFm/qvJXzndwdhvpeuMLHJ3Ke2HVi7+ag8vnUF2+ZQEa3gbBiOAfr3J0Acn0+3VoSDwYkE
BCSq4xAUN2yjAuqrGmFI5BKcl5+8YIMBnzmzH5ixSTxrmjs+qCJLL/w6K8QtawcRKO0XalPYuSC2
gcdzECerK6LdxwCPvJdptENkPhnGDLoG0pCnQjhflUxbq3xGjX5/FbuLlyCTuPDDl9i32qHGdg8B
HsK8vVXifFjavVQfrHYiy7n67zE8VohuPph66+sr+VojNxwcCCIRa8KVdWy/S/3wsbGMiMs43ZfG
yVMiS/v0ktazlooECwbnZGdNchx0yp8/+52galGoCZbtGv09DAQlrtiDj5wMK300KWq6M5406EXG
pyoeGkXkTV/2BOIxN7r6Y+9+6VjizQpNqdsHlrECe+PIwyA+TXGE1vQfxdFAgAZbQb7fdxGrdWc2
EvnHaEtKrUcegye8aZLAtdTAlvTWKkVpVzzUeJYe+FELwwHfRrQ9Cs/URHQdxObFNE0XzNi4o23V
r5Cl6CIYaErfdYDNV8Q9nri715SKdeXmnOhNyRPxqCXVj9NeWfZeYcxeEGZjnIqn7vTP7Ef03V8m
cLlphYinmucyZKqyMV5BAuFIVbnA1pYm6UPL0naQJ7/CgVzFlRDLeg/5b2oIw7GjBO82O+F9SaB9
KQ2iGFMOayjNcX+JptnnQ3QEdONFC83jSO/4UK9dHOC4lEjBgqq8svtAJWG9aDKTi8jiTvvsgWww
L7fdzOq/AtJaNms+i75crbaoQ7yitgeTMOkWYnOrQBYCG7QBPTeabc1foKA0QBDW8aRh3WjMpmJW
U5E5L7ZfDHpZXREoF5VP6fzzhzjfz/vkD/kEVwEF6SMAzohtA86y1jGGkC3IELh9nv1as9PDjoh1
rNDLHTffk/O6CXcTc6Fe6OP0UCF1J+C41m3ExRp1P5+/+k6B6TxVzrk0eAw0E8RO7k3P419dGci7
zZNx0dRzoCVSnphmd1uNPZGWiiUlWyBgoZUks78sEePbklBCFe4o1YbeB5DhoB6cqO/9h2raKhtT
063tdOGG0+oQ/9wc2Me1q+Jlqy+DZBWb04E4OqLQpC+ZFpyZnvlxh+A88JfU2ETuPeW+fw6GZ25z
5OWUYkxBRGoqDjB5HUZ+8gikpp7xtSHHnYYniibRDadziQv4kYtu/iz9Kqa4L7t9p7Y3hzJRqwRy
7rSOmKxh186x7kW9iAk9QwsS8oSJZMdbPBldxn2pmqG7Gvt3m+ZwCz4Mb46GZDW690ERhCddPHA4
xsiRx5CZkzQmLSHoXc2EO3HUNsCJNPCZ4nNXX0NWSgiejtxknSRVvTAa3zMS7BWDWxooOhy2QaOE
EhAgaFwh/aCxkvFxky5XJtD5LJwetohRFR02SaYT9IAI3g7AYNauSsMwQPK3CsW2FmgKJsxRU39E
waVPgP7X6CE3gdYNcBoo7Ni9Ny49WT+X42G83Q8DzQuphO4Gldl/W+/itvYNFHnPTSCajDTbK2j/
z/4On3myDdUz5McCiKY9kabfsubfMSfxZCM6iesd/4kyNGkLmAM/7VH8Ha7nXlutUOuzvh34HMIK
yMlXVwE+elbDyNdTAwSGNNA3DaOP+favB6hqMSxjYth02Rr9BDLHy1m9HL1UBmvmEIH4pjg9lwUq
KwkMKiXnxnRoV2ZI/ulMvzDBCr/p1eaDw0ABY0YkqH5PAgH7A0EGqfWq30bYT1kZGn0eQdkdmjmd
TNLHIxHjgWEklW+MNYEj5zzLDbVqtdJr6wk04QkW4ivxtYnzOOnRnVXgpQoy3utIJqigPwjfLLp+
Kw6NcZlIbTsXzyDXVKP7GUc47AnKB8gaxl5VhqzCa8TsCGfC/KMgAw6zzGxgeJOHfOwzfsF7Uoyl
uvMDLDoVmarLsQKyCj8CH6CrmTZf1NIyYKBxf3dcoY7SaENjDZSMFdbJlgfNlBmbAdlpvdZfKVcS
VcDqxLo7zcVkcItfnQ4uYz2QrNIY6CXblmcd3DX1w5AkWv/PIQvmFmUMdz2/YgqDEQlePZ/sLd1h
0xB5NYEUEwapA8i4ZU7G1MHT/eFoEoFPYOsqLNZ8+OV6isCmL1Oydmt4Noa/yVSMu6kGSTvabfp5
C1Am+UPczkEta7vrGhjX+iZNuaYHrmrz1ynXV0S93fCwFIu10NRs2aad+T/LIzwI+qQXy710/lWJ
QprzE+FRwtLyXySb8wqIPFiIhIMj6giNkriFALaji+OB4xTFQMphWMFCHkusgN+scxpCBEznc8M7
mmszPApw5wBgO+2YIvcPBPi5Qn32Lk8VGjNnPUuMcBCecApy8TlsgZ0uNwTXjrPAq9Ow/3zHKjrj
SkP40xmiZWPUW7+zaWTmhaT2bPqqdgDrFLkvvVc+joxsmzit+mlfe/jW+d3dLYmQSVOOwBrIHVIU
5V42pZv4h1K+VzsXTubQppHWE0QVwAkN3B1/LUz8GxXrqNsoly90SR0D827Sw7g2lONzuG2dD17c
YOEpgsy24zKy32A+iucziAU6W+2ulbTidv3rlislKb9LZj+VOys5BCoON0Y7ptfakuSl0blv3Bmm
wGeE7aCKnFxjvoT5WUnM0ab74oNJLljw4qOaftNN6QyKVnyWo53gr8Z0M+aw4Fa15gw71RZwbXhV
RtEMhWytEr45DfO52JAR1g/k8JD8mqgJb4NmUgJ+vmgLvfzZVtEQwxo2AEaFXv8a0W1WLLsh+JBk
VvKzIqu1rZ3hybfOyWa37WIkotZokXEqwPPjIY/KwPBTyeKfCIsdAs7gizF/hxhHGHy2raQL8HWv
IbI1wTZ0xiLhvWJRgLpKAHUIxhrjQX10fgUroIgmrOWtQHrielDkZuNXt6e+PQtyt7eJ22g2YlO+
rlyKUrxkafNo3snK33VeRaChwLgFDqa6rk5ORcXjEnQfT5WMn3sV1Unau1SmdfHNS9E98jv1s1V+
7RyMcutDrSwag0h243LrcuiVvK+gjqju3CX7ISj4h0SG+Q4Exi/iQEbMFcfu9/WZRKCBDlpEoNg3
qm5LYldZR+keA+AwO2reTkiAJ52uCGENKbdTwtbqg0SWaGQpu15khQbHob/qW1JB2UNUyxHHBkoN
SsdMB8z6V5Ta6N0hOyiyoRf6kO9ubs8FnOvi9oVZDSAM6gPFNFrk9iOG8YChemlW8s2uMBOkmIJP
Y5nOQ9IGF07i27iA/ss1Miauxvk/6Yd6QfcO6OTcFdF86LkmZjYngLD9clXqvrRUIc16kOBzujVQ
vBYfQ97RaIFE46SIf+U2WgKHAcx4hFXAtUERwQUYf7XmvqFx85cwrDc5q6pU1p7w/m7yw2G9Im+X
2pCLs0K8/zEhNPy95XfYUn5/H/vzKOZpKgkgz5Vgf4/hkNI2BjXEUE58IIKa+d9HvFEw1HeRri4M
6fxUIaIvQNYBqR0bQnRABtGjh1LDBXH0naGVXy0Oi9ZRt7QeSqcFhI0psmQQ516/IIpjSpwUYqhl
ugoSzHZSWj9CUo3T5MHOeiXo7kN9gCBnvHC3hsaqAnQghBK1uGF2bL7/qQq9pknoj1QiQUwDQ2JK
56/MYleL5U/h1Xlx4xoAL6eUV8+I78O3cyDU61B5fyXGsd+hMOymT9YsK5/qqCJpc9je9sUWWMsk
x/wheIF/wzSjfk1JPlA/VqV9ajkYszALKCsr11TsKDJ4GsOBF6Nfo1PEbtzxpfunSZUYRu3SJMlS
brnu/e1fScdfAbAIU+wJk6/jg0OZd2D52qQ/9qxr144oUGb81pcaqCiWqdWifgR1LZpjASLPnTZ/
pYZkJSZL53EWeTtsxj2NRpJnTiS/b+wpDF5t1ePcEgxOn3H6AJManyGT1j55NqE3/KK7eamEMuBo
EILA2qV3uNLq9XvfZ4Dx6ILv6RokiGtCnz3AOMjqWyJvw5hVFho+MN9WFzYAgcrQpJ5xV9GUv56g
yI3gLpF6H0BFKbME5q4214N3pFdC2FiiMBOB/jPuesGpxIRY2/nyxzxL/d5jq8+yDpyTYeMvRdVd
6+X8nmLOIvxYyg+i7V3wbA1V3UXZ4jymAb5ItAQQCVwi+HdR1QMVppiNOLRigO71Aps/mQLbro7/
SuMSQeyoe8DkHSZWO1ZBuxZNErs36Hs0kontOEOh3FeRTO5+8WlUHTqkzZxWKnGB0Tfdx4+qCvpf
bAYluVpIgXVYmWrQ39209QObn+Kf/JEZowyj3r+lUyw1E+k8tKO/4bJOQofUe0U4oQwAXa8hl3WW
eXavmR7Qv42CHGU5BO4mvuJPS+/CNCwwo34aUqmcNsu8PMJ12wfIzwBNFXP+BL3/pI2VYCwmEtOp
3I5dNjBwcZ1LLG4vHFK4I/oZEMItp9+kP2+YHm067UVcFt8wY8hljtViCzJ8oM5tQ1O5hZUcLlyQ
zOMlnPSPZTC4pag2YtlxWIulvqNsG6lF00gOfR5xQRfYECy9lfeEl64Gtpn8S962lRCpid7ZAHLE
47HCUXzlr/iGI0QlUTvltbSBCTXoM35veiKZ+QrmrGqbpaMyKJ3WmrwGrOq5B0vduJAOqj27yEzn
TlIl4h+PqQTZsDU1Ae26PfZR2xKy8ItFfaIOz5Cje0vvdiP0sLhQumBnvzPWUXRROgkve8CP7ECb
RtYBzodxs/c/ZePR5tDJarq6IIjiW6TDb+UzMzZbF7KFv6Du/atUysSoob0JZl3pUjP526b4bdHt
ov/xw2frkq071H88v6ewsr67dEaYnEhhB1C1EMvVoovyKd8k93dZGQsVsiVB3dV7AxNQKtWqDEgb
EV5WBKTMZ3yeSIcwphjKOPp/2U1JEcX7ylly7zAQfwGlAgmY8XK4z97+yWJoQtRId1CxmdM6htor
iHYSuhQZegUYnjxwMSYRUNAtJdzbyPNJkq2cxgzttQdoatTj7Fkkix/4/8gElN9wS1Xmlc1rK6J8
TOJ6vf73y/B0+0AQrmRbOZhhL5Ogp8vVO1HBL2R6fF48NZVXFh8+pDRzUAcoHpaUtHdOAG/JO0eZ
SuMHuMv7jPOzMHrZ0gKWciPH0L7CSjrYXiXUsI/+J499A/SW3kwBo8PiKLr7lCVkJ+7RX9kxnX/k
0ca3zMSva1zC4gCVSXX/lduUSDzlaJINzL9VOOkNf55f0fDL4vHgdhJZlQ8PB4fMyjlpXPqOdIRU
FV+uDXCaKvAkBt4HgGj6h/wLbL0cvBqM0FR3i4bagWqHkFC8t6QEwBUFIEKAkHJNtret2KZxq1YZ
HUSl9/CTbH7aNvPw8fCx0q13GzY0cdTErsU0l3MOV4mqDq9+7e+4ildYQWENVunH+d9Hr6deY/yr
B3FexOd7BkfxveF+0/j0zybVMi1bX0yp44fRB4QLU9Bqj6NdTz5Vd9R0K3tjev1pbFUV2PHusFIQ
5pCdtW86pqEn+T1Hk2sUzmU/Ea3Rm43dBQl43N5Uh2m2YQllTeZVsZaZH5NVNG19b8WKg7dRda1i
MdI5tFrt0FE7OKuf4UOU9rsjljygtZNy2ylHnsw16hDL0VpS+tLDdVeU+1Ya8bhgBUCyhVOFjNiF
bcGKSKFbwZxsT0ncBhuNINxTrr5d8I7K76TEMsNyBoE9OiKPq5A0aa+4PcpfUZ7Pf26jqMMPYVJZ
3KpOWZfYtzJZVmEaXrMCRAcNq5e0KjdbydJqjeKq7a9v0sGkatPR6MnZUe4OJmmoULEw5ZxnwjFW
WzZtK14VkOfPEHskMk6/47skjEL2UxTDLV3J0q20I7EW2DtMTRGnT81E7xeSRKAw+uUI2XMgOcHc
77XT73cKbnPivaR81ajP2D6XMtOAwuAialLlDlHgnFPf5bi+J+a5TmMLxiwfWeaooTYJcnFVdhdd
r5/jpLacFHKAraPIHj5GRF2buGaLIlL1JpCYl4NR9mcK+CLNr1sK2fktxU+992F6raJRdbv27uLl
XGo4KLlDgt0Nc1q9rubWni22AoN/eWioKe3N7XzPYZnG66P7RTJsOo9xWKFSQDUL+ABWI8Gtk/F7
pcZmePTlaqbFR41SiAFcI2wmi5JZBGMJ+zk+YsvY9bF5m+P5Lof/xxBffl5CDBTKQoigGWcrbcoO
Y+old6Wu9SvheEDqAdpE56kPjdaPauW477dTvwesEyBAzQnODQNasKN/vqJlNF360DWZfKBCCrn+
9HWb+RWZZE/Mc10yf2Vwo8b4xsbmyOGv1/irGnFl5/dr1e3k/o6xkrAkqnOfCWZKwv2jmpoRxcbI
Od/ndChmPPcr30L7OXJ1i+DC1NCZRG79+FUVEDqt/0DfC0nk5LVALFL8aIqdpgBar0LCGGBpH7M0
gwQ1m1oSTNtbDwv766OozhVllA65bFPhO/I3ziU3BeyM1Dcl+HGNtkVkhV2xC55aY65H+gMNIHrn
x7iEObmyo3wD2qXRFwf3UsGAvUZ1IqjTRGUi757VSVgrVP/ClJjVWWvxx4/GKhItbC8HURzaqFp8
wZRsG19G9Dx+OUHbmKnISxOM5EiLWr56D/jsf0c2WYrP2ZjsIbTjjsGNCpHlabsxNRxnoC2fvkgP
lRdJLgVFOICTWZVGVFD2mjXyhYaliLltlv13pdZZrKDHusVb+gUpByhAnCnz7Ua8NSNRw3Zeof+U
VziEOfdLVpLqGkAFCZmtdcl2t7VJHu0PWQFMOgMAxAxs6rqGY6+my742ZBdoUl7200YJq/MesxE0
iyOh+aaAjv/B5sTTwHXAwwDfaU4YNlvm8Yy1sBTCTBCu4iNgFTe77uKgsB59/gHxnBi4hL38zj2O
wCNfKZv7BZ7sKIi/IVFvgJ7bNpZKHPENRyX0VHgnDU+bTf49/burGKGn7Ok+wVrmqST7jK0RsmeQ
uYY+rWF/cZE9ozGsfDNTg032nsv2EKvyUn5yYQDM3WRlOgfv0T0tXUfSkuBl6hEuHftR5C/YxE0D
ZViLpnUR6sviGc1ehxCsvVkMzqnVwTccx4mO1LjEVhRchGZGvd+xeLbqlRPfvs17ELuXaDOeDyt1
hMKbNmjt3Wm9N0nRzMVsuDizbrZAVTd5huzTU4FjgGKr1wHOi57klCMrF4U/RbgRP6c7JqKeM3Lh
oPU0T5VA5iARZm+603ydBJhh4x8Y3439jstMs9yd14YYctOpWaPfUFw2aSyRR/mdr8fNc4cMofgN
ENO07wZ9USAViSFRyX53ln0dYO4N0iGbpmWccArWZp71sZfRGpdVJ0qSwXA+kf/zRQi5RcTvKI17
Uev7EQJGdeg5E3Lde9VQXfD2pXLpPzh752euYEbYpQwDOFnzjXwL/Ksxp6jnhj3BTBa7Dz9kSD/F
AqbT8weDbvqHo7qRmgp0ePDlA3XjJCJmkNcOQaBeRkfpwElPEA8j7cb8xP7q98LlAthmYOmySG5C
szcNFrBUEvUBtKiskD1uCWu5z6nZ3u+9SL6NbbdjIjxgpONsdtPKe+9q/fFPnhyAbam5iLkyc+2s
0zJkXu4mZN1T+0Z0sZjhlcS56s5BZbLbjMc8TxOBySLryNS99/6tRg664SP32WoJmZH8Ly2TGKyZ
5vxBl915quD7+IY2MareB9+xdvgbEgiTzslaC0LV1MIA+vmSCtz1DNof79KwuABEA3wyFngZm7vY
jC+qKgXtoMuwBzOYjLbuBSIjThJEfm3nWJ4zrl1pSigazt23i3F2HtYAtdNTJkQqlqOEQUhKU5MD
bp4mT6q9VpqGnQsPPQCR1+3m0X5dLR2jQy77noboi2Aw4skfichs4woHsI/thWdi+bjLx9x+axBh
0PWAMsrb8DOQYCFlvdjzLLLTMf77GGf9WhwuA42LNUWeoh7Q6XDjGzOhPpvgwFPb899BMZjNo2hb
MNoCtQYCrLW9Pn3tQTR1wH50zaP4AzdE1vIdjBwPMDjIwjrxQxsLsXan1V66uiSWtdqaw7phTHDv
sl2Lx8GFYWYvMbp3bwgYLcEq22TCSLN02qE6QQjeOA+ESdzMm1C0i0VfrhRNrnhsXDws4QK9kIsi
BsQcypscUafhOrAPG3Bp9LXjcXeGyBaazhehz9RuBYHPr5bqJG3v5rr16JVGSjQtxSawJgUK097l
jo3fxE8WD8LDHhf9iS0t/UCJwn6y70CN+kdRt9Orrf/AwGiUW+LA95Nfmxb6FA/69WaG5tYz585I
UOVK34DcIyW44TPQ3+HN/nDOJ7i8MM9TnoKmJiqvq8WXrCtqy18jdWsv2nmy7P4sCCmjM8mIuxOD
hk9W1wpuaLNoKjZwCEcQyin25VBvCcNKHmvI+qKGYyae7Wj+ORx8qsJG1q2ZStUhuO1mR+k0YQKC
dHgNEdXzT2WkzmcGzoOfmLtlxnIvo8vPStsq01FgU+2PeL15cnQs0J+M3RNnby9bHY3Ti8e7BNU2
dkpIPseBoZAA1UvmhMgZUEcegSafXLmoK63IcY2N3VUoe+WZaV48tf7JfVCZSnWOi9+n7yx0yKKF
HED4M8q59JnToUqtzfTOAX6ICTOhhLCIUYWKU2AJjr+7M+PqK80Rj5fDXT0SoOMh2dFuldc81b45
fZ4Kg2cZjLarb9+IcFUKkLPqmEf1QxpkQjAEFaRW+pphSjlhIAiC/ShB7Euu9gbuuaa1BKu3L7LY
o19VAyRIpnc4qUiXN/k07o82uaULcq/BR3sXx9QEShGFIG1DCH7flNn6Th8jOc4V6Et1amHI4PPa
qeqaKLkq7ODckHQIcVVCPAo3kMZoUp/4fDnIJq346rBBQ2KI7YbZhYkQ3LTDX8y1yIaZvLTANeeH
2IvrtIQFfAsrLBSkf4W7DzE6DFwI0D8T6uEV0G5lJHSowvfq75M65ebwq5D7ijnRB3fLYWrZx7Sc
5oQIHW6BFTJ6YSUgIqVLnkzrM8c1ssxocAFih3HOQWOc7K5EBaEDK4XrRLjqV8kxFrixywv2ezna
3FB6xAb0d8RsBFp6nXst/fmYBxifrBF/hBrvorYaWnt9QTusJjhpTdm54AcVGijtzj2hp1+aDqAN
l7k/5IZRg/Tey22292qTPp69bQOcxvxNBXbD6l5J4On61jOq3bl/KzwJNjCiTXLOvrBz+BqAqGmh
THvWgacj5OCa5V8A9qzMFFPgCXB61AGHMYKjnPE8O0ah+HFT6nSOl7GcnV25FRofFzVyTTBz6FV7
epgXJh5eZep4YNX5EH0v+gS+BOAFPEWVdzAlg6vG5wb9TTRFQxT2ZmT2SM7PILLA1uaa52nv5K1N
xt9HKoy/yJIe3r5W3D0DDvxohMrKt31ntw/80ZkAloO3OyZKDjFQb1AHVrQeTGhxaxmcCnVisy8t
ky/HzUOuv34D66yQcLr7MgjQFe8erysQ0O30SW3rcUPWfHVCv1zqTZ+OSTqSGgGMksKXCj/Ndopl
kBKY0P5qwlyqYfPK/KpV1xogaYi5Xa6GzRtmQVQ1MRuJYijnO72SsAvPVHgxhfJdmU6eOorDqPQ8
6Bx5/LbOD8Paw1tNOhRMZPaTcp52eWL6r6OQ2xwszNt7s6KOMWM7wG8aStgcrzbwLxn7DID/we5n
9EqcVxUz3uM+o/huluTh/6MivV9MNKfktz0LltxGcOdV5vYehmIaK8r9MFjoiwM3K/DfE68G5Hnt
B4mqLZCBtMPny8SQyVyJfIUluX1VCylFrHIXGJPsgpORrMjGKpkSTg+iwfRsofcokUt2tTMyvG/h
iKqBu4XXVBZm0E7AolUD/kFjWyl8n9aXbHPc4J0s/cslzQigHR86TP2f5/s3u0+lrR0q5BFVWdC7
EsPJobfVc+KbmnjIk/95ZKyKbvRaKX7BBNL7pS30uj5fk7gmpZ6S88B3E9vK0ksPCTAwEO86MPl2
u6NM4z9GEUXh5M7jBn2iQzvn+JPb9JIOv7wUkvqcO1BV05hnKjorWOjgwwp6ECz3yIBAA6p+SbI9
RmEYniTDqWnNVczMSC63EEGvRN88rFGg/+WZZQTJu6qwVJyE/kw+FeyEoudUMCmoXAgMz3LV0mGw
UktdzDa3CgAclXUNgznJrQUY6sAl06aR0BkBo+PBkENsaP3sVVjhZVHM8hZtIsv20ORhklmUqV4L
bZIVGuVy88WU0lQLvIPjmzVgXJz+TYUhP4He4uIB/RsZnBHmQYCnQyspHOCeY9BhyC9dNZNusB7d
pv1+leL0WzhOU9eV47n8KyE2vlnQEz3Poe/ayXx9AeqoaAHQYqmt0n4/LIydUDeTFuth6WC7TSSl
EitJy3gEHVzPDeoW84pjDJ92/rZG6zMAAWPzxrOhAh71dgrRWERmteHcMCZ/Q4Do21v8pahl/+l8
UbVt1LSCz7lcINhtobUB4djYaa1+9fQcp/sGbCAJokfJtNiX9ys09BAaHrHYJlyaM5wmPrKd1mq/
lPLuo2G1OypFVKz81pCxDHBgGXBZ/COmsLdi0kF9SZ13rZWnz6T4LtdO5qm99i41uHDytWFgNo6R
zyK/okdXdwAa90hSbZwgbbfBZ5ze9t8bNYJaZ9c78G7gKtTyse97wzDf3YBucXh7wv8UpsAZEtrf
1oS0TY4fMiJQ1gcje7DC3HwQeKPPTp3ajjFiMGyB306MePw6ndRmGg1RzYvqCHJzJUFuUZJ6VPol
63pa5SD2BzE5ZyT7L/N8wU5rjqrNZ5LxwS2zmK49NmbssPF50uydGlFcW8DgnFmkDwfgI8G1NaPN
kE2Zli02qPPH9z+6KgqOQ9WENg/Vj/xATElpXYFMG5iZD3nld7iTlA3dsUlZMPSZrsNPn87Vi/pP
Q0ZwnCxD4FhUddKntBE7ILp1IsBHRGn+fIWtObXN6NdqF5Ke0m7iICGMoYaweZzU35TqhUXPq1DI
7HsyDg44eijbiojsA+Cbl/sDIC7xA1qCQ7BvnvRyg2oOR1B0YHRF1B8UDwmGy72Mj0L0x0+lccJ4
kju+9eQ22nOQ8oOVJgSdG8FI2NlSjuwQDvtwvog1vQBR0dpHnGG2SafMCTxw4ja0jOHWZMzOUatn
4nCfacvqPXbnbzrp1hF33ey+a4SPQ37td1/0CiW7zt8jYgUlz8htbqfBzYZ42hvJ+ELRafSVfz66
t7ABacIuaQSNXIfX1RGubnRchoj7zOCBWWkbuusw1uaPmBtsA8JBQkWwpZye8MGxb25EeU2MN8ZA
8pAAaRHzWGrksk+hB40uIpFj2upWaQ8pI+EcRrXTcfgNpSqi6QqZ9haXe8lTZ9KRsJQyikFGuvU5
ZKleL/pyq8kEfJQX5tLLV52chVUO+YLTNEZE14Pcc9swLf5tY9EZqAXzVP8gNCCU9BNkaljlW80A
snulsLKsu9+MbGdrP2K9Wy/KRSTVt0Ss3MPJh3QbsZ2KzI6+TN29puGVw365XIW/l4m/tHS1IeK5
Ch3xvNvD+C1ddNDXF958Dd86HgFiwYl0AAOWL7fFTcfcFVMUL0K4yuBTF0jjBZhuJ0Rmw2jW7gg5
c2nL9ZWnQTBa+t+AwIWYGYkD2aMmItnFGA3V5DnvmofPNpodjGHriW7u140+3A6pElG06HO4fB2e
DjJC7QtbRkzZvizN1sWsoL7qRX8O2z5huJOpti2bSzS2qIyh/tJYbeP/lWLZ7RyVmgp1v4QJ/WWl
GlWuhkJ9WxGOX9WBRHkx+1fuHZEzQL5Z4oY0y8DrgTILAEo675h0Z6l5/29942bENFEssM7xjugp
bH61QlwR8zCX6KXgxkQNWrtCE23pVm2Ud8/93d2glYCK3y+ctR8OR6MXj/ZQsYK74CSbYp8yf+Zg
3BYPhQlI009bCoZZUeQWmAI/zn8NzikuUFz5ThSx+Yu3r8b7FcLx4yFXDcLigegquCR3rZZKee68
tQzjYaV/k3lgc2ZPNdEQv150Ny63cxcA8jq2iYcKmoESLRg56ZvYq/9g8RJrUAVGL5kBDCLsfxTW
sF99esZOVuEKP0lgG0gfOkt7fyvNS1j/Lw+rVh/NMXo0NLKxG06CKyMG82XvxLLUhINS19YKtltz
YuPEhmNXFRchLl72TB3DL9qJ+G0JKTV1MRicf+dUFKgOPTKGn1Key04doWjkIYU5zzjpEKXQD0R4
f4urNl8goTWhcIkNE5wuE5XGFEbTlgAt/xTzAjC8al6wMhGefcR8znRuooGJhtzlI1GGnUCV19U2
jHI+a1Ii01YCrrQ+cRxaVhtunHKBPbbYU0FCsi0jbjMngx84+oQxjKesm3ojkuxv8bT0ZR+Azoza
SvO2P55ELyRON/YhSTOmyIFw0wEHgLijFoPCTQga9X6DuZAyt4pzo3b5v199ZHmCe3kwDEkP3qQB
WGwqCFCA8934pwz5p05iTAER7jVmHFPjwVqDR93+bIJxg1iMMR+ETKtrnnuulnGwB/gACPVdnfcR
DiOiKRtQW+SeU+cxYGht4Wwz/QCfE9zfyLRIfE18+cfLROvBbdrO5iXjLVfi2w5sZr6F7nCNSzoR
BTm4byvxasN4bxqZG/hdP2x0jIfGqOAeZn7tDPs5ruwbZaJ5JKX68TBvKGxJKggdDIPHN30aOrvF
gP/UwyixOvIrzPZnCdFy0g0+a6J3qBWqgKq11gMa3mqA+rWoyX3+lj4lClXoj2pMQFvVsHU44Scg
XCGReSfk0wf15xENQX5dC4Y8GjNiESCoNYVpwK9/pMhXcCoQk8bqiqJ8hor5vKIDbBhjpgXiWADc
h+vTlu/8vtBOhg/7z4Q4YkTjFv6aLrOAi2af2dcIqz8NnaHWWzMXGFWvCETw/6hCwkApnFECi+sS
yJ4gC3wH+QNzfvd1qdusSdHwUdvMFXjS7g78mT9pUl5tgtSEkMIM8LEMYkk+zRrlfziaTN5tnxU2
K/dv3LxmLbdLmMvZbwW1q/7RaTEg5EM7V+WkeIzkp4vzP4sysR0Z8+5jwHydtGA4JaBEeCoHa2ga
9BzzMEOTFfhEEeW4kjTthINpOL3HjAo/vSsNK8XWRijTmA4DkN0ZCPXSXnWnlHu95IoRo9bJOvkE
A1+iBOrxE5aEb/yljNmSCJtjRVy1wn1gGQTKFYrI/MCf0lifB9bg3P7exL5rH41KPX/tcKHpjAz0
pqO7m4Ip+oo/W/24pzfVW+50hcylykE4aPppuodPBkFyF8uEYoohEg0UUUtRBZgUdubOJKR6b3qB
YHuTlm6utqaqcihlf/CWQxTsWeD0njLlRM6fB0dWmXyBaRzKJ0IiQlTX0kzT8EJ9dpNaM7PE7Qqb
eQj+9gzxDJ/8d3UUiOoAeUV+0lh9d2y+TxtE+DCtSy2CHNBwpc47HpVkB7TNMTATGIABsVWYifyy
llv2kW8ASLrZD6im43zUjvJxaWrYApJSz02TzTNwXg715WSNcildqUt5Zskkg1cW7xMXceIrY2WP
gkyDspmGJiqPX+qmzT1fUc50rvNRceme9kkzn8DzFjtIdfzXjh9wRI1jYjs/I0zr/7ofmcN74axr
/spb8jP+jCJPIg4FZ9seBrYQrC0PHjJeqeqjZXJBYlBaOH2r3N/BkO8qkNSwQXwEmSFHLEzaLr8b
B2s1d79ckohGuSJPtw92YYhtYTH3XBGbeh1kGVHKPAN4pWhCXBZa+YHiW0lo2jujsMRw/PjdPPGP
RgQQQzVj3zz12z/4WEg6vesrdhlgyRHjgA8+1eLnlppyuLdqtuFW1+5SeYDgqnAzz00SgOtaYpIk
ODtbw+cj4hGvKIidfVTqymbIQeOKJZlY5t3Y9q7jftpBQkhDH6MvG+6mdg1MxgMRdIhYTWB541lw
M3r2U7AyoT37ramEqRwECbkIJm2wzS7mxOWqRhIJ6say1fBW/EoErNvwD4INP6VM572whxKL2UTt
DVjHVDomonapNqBLm/v0v00QE2rkH93hxsHWD6TrvYPlP1iHSBhSXYFDcjz69uLIFOiiisNZ4iV5
BpYMHvdl7JbrnDzDS50mrkfRMt+1ZYhDzfYK+qt35Pbr2PifQFp3zNovAlLfPikFd5Eil39ORctB
GjoAaRDw62BuoqbzaAq16WoksCNZ+43D+fkJpoGUa3jF5C1IT6CDqVn4CzkhTYQ71zlv3PF4lqI8
Y3YK/VcjpY/5U+vXrgozK7aR/UkGO5yx3VWOtNAOBMomeXU3UYBTtaQJ79QE+A34Uo8ptXIejlHO
WVwCibFztQKlj7AXTSo7uBhhk5BrIRKp+zM6BelC1kNHjMJoGJQc//zVskmTJpJ6hStzymWwMZc4
9ihiTwFiLAKMI7b8SrlrQ0wp8aNuy0h/AyZ31aB6ZzX6HJ6I3/bfP6ba8U6zLrnup9Sgj21l+Cat
dcHwTGIh+TefEl08WfUD1aX3tdX8YxuYPA33Z4Y0TLiukFk+zCIfUCIozadJ+12MHHezVcTPkvPs
BtlCcb/wSYQWXJsym4kV11G+nMPkw4sp4x5sweFh75O5UACkS9pFp+oCtbUY70fLgNAxBfxzvVjV
dPccPuxHKN9I9htOSiebHDanQorZpZhUJQs5S9+hX6fPsifQRYkcKZZNUUkd9O3WE3ny+HQnBukg
AcPwLony7lvsZPzuT2oa3GgQLg4AhqbNnFidUYOSi0g9SbjapsFrhjf6hvDxURJQ2u0+OZTj1+Ho
xMGBaorOILZZXdOW+MP4MV8WdoKKz+EQK04TULn37zaaoxyJkPl0Gbv/iHWBlJzk2PdbtxJiB9zI
Ld0nfprULFf/uzkr1TyN7jGDH5nVmoATk1XJ207qkFYYCvHY3Lp6CDoma/JwBKWfYJc6xNbmQ0cp
QM1raeail6pu45zcVmIwUh1YoUZyRF04oHtl3BuG/eCAaycLWje2ic1fDzahh6dwCCRHhH52z64P
t2x0rcix+9xL5u8hnrdX8lqIs7/ymUKDknVvlFW7SbNqf36coUIBrmORpI4alB+9SoSU1fCLL3Wu
qnBKBch72UjcPBFWbGRsdKlU/+vSzhuLlFieenilaqTXPti4PRIblfrJ+sEP2ti4cDomH0KCsCZc
vXT9mZQlFFKaDv35Jg7onD3Uqv81VHzl6uS1phfiww/D6Cl8lbLAfVTmVNLcDlyZna3Da58JZOx7
lJyNqprRXLkRJZaK/mPSnDcfhkQ0lJ1Fo5ZguieDwjJLx4/lPWQRW85L1WrEEyq6n4WQdvwLFiK5
00zqL0DJz4LijRbleBdgV/zJQJQTHvQ9hbJhOs3b6cyCgCrH876HO8/sIQAqkhfg+MOIjW/eUZP7
wycsBjooAVM6vfCfEBAPSV5XofovzN+qtr5YDQu+gy3OW81U4DvSa/asUZMcxfi1s/PNdLv9X/8w
hNDO+UDdo92I1nOEPvasF15aklkH+JQlXwzQ/gQXbE6Khdpt8IbaakV7IDIIbH3y9E4ww2A5egjr
W7gocQD2TAL2e1vxaKXK4iYCRv2H0PcOUxX4bHNE/uxeHFe/o1elAamqlGge4CuDQ1rufhTVS9Im
jbCxqIFxRGoM4dLhF125pydtwgqZco4CRCIpJDGmCJ2MGtR5oAcgLIJCa5YexKoad1PdHnWckDxV
647DJOHG2J61apjCF3fvpi+7nM18HChpSpdfXH9DMuC57fa0190ttZ8Xc/e8MxOVKV2Zo+dlGJ1w
+MeM9INN2aVp0Ir6vBtujdJdmKtcNnQpjEWvQm4ivE/SRO+7x8zxcgG2xFJXVnpHuo+Ny2+IQheD
aM3sb+LEyjtkuDLSAIksdW70q7EYT6xkU3RZ2nWEsj7pfj7BSIwzKsWMgM3xpI3sAlIeoqFXWIZj
JsC2GpkxzlXCsyCVBZ9cd2T9ED9fjTCly78ny0ycyM/VAMyOZzILfxNyDb4O3QYJpKu6FW9kQbBz
SDmDsMOgu2gjrb1neK0MZRioBhglMnGg7GpJO6+HCJFFfEdtVTpUwlxlojBkjHiQnZPZEtk2onar
N30AhvIvU/Hsb0BSK1iHcVTA/3rEolbjXS0VK9p8E5yr/0SC3YRX5tWT/NHQ0M1n2G8VwmG0oGn/
mrAjEtd/E7g8qvW5SgdT4NLlCXeK0drq5/xvVGImB1sGvUsKMDsKNTNPsin2Ixvx65SvXOYncNFR
cGsHCusz0hjNriQkD4Pj3xCEuwQPJ2R9S7z1qw5TH6ig/e+M9weDuPfMf+ipmI+mJYgYFH1VRm6L
oy+chC2xbRqUtg6FlvfFIghGBzZpIGHCH/Qo29tfV8Jc2K92Z/3wJ5pgV2aa6IqayzD+U06adHL+
EWEvzOf+MnvsYCIyLVabQy5g5Su3DMVgEIVT/MlAlTEl9rjD4TyTO9nK/LewCfgKFaJGli3l0H/o
zVjW8HNTATC7xUQ0AWBtyG6D5QeQsLIRbk0utUjPze0ohBOnYp1lKtv6c61XLse01Vh6ewQTj6xo
nGubRhgXC+mRb4rR6qWrQrdNZWRQo3vf4r1Sq+M+c8DjQIfDct4fh73rfkn5SIoxvayhUSOoBv9z
gMmT3Oky8A6I2yh6rq0iyoLxT7OmEGy/Ecraltkck8GmyUDOrgyW1nPEQnyWPXoTIi6ZiiCbQr4X
W/JRTAz5wwspIRpBiLnaOYlL+5g6ALuwBX2GjkuWF+PflgH0ch5nWvB01jc2X85FyYQgcY9OCBhO
erNuJfK4sJ9dy+RtlnTZoJIZm03Q9HYGcZzagsBFWDtpLR9BrQQ1n+w8z3cAuWxmZi0N6k93bis6
miihIWYUsz1oA7qvi9iQpg7GQPMWjQquZOugcsKt+bOCANHQvWs1oiYP47PWrAScOVZtJL5gzS63
IsU8XAVjnXS6tQHQH6FW20QO13M2p43qrh/K8ZH//Q0P259YFxiXNRrfFvdK7GweF6zJRILNnc6k
99AcfHUZdvfXGO5Ci5W5nufl9PHw6FzWa86dg+paPoLJZUFEgLtoE2z3GxbmrqR1j2fJDTDTds68
dccqlNARx/VwqwA67mSt/A012qMgP6WX3rtDcoJfyBhpTJsVdSpl0GS/PGlSCXfFUeRgXEKV7k+P
hzorBDWFQcmeFDa0MUc0KzwLP1HpIi5sHND1e822G//mdbdM+xXB03oWr1WCfHmYA0iSUsV9Tzh/
qe/i4DRc12QR8vkn3yBkIWNsrdYQ3vkKwJFOBT6Oy32B2IpdTpZixSioAJ5TTrWbkcZfyaQBtanW
uqBoiC+UM8/CedB94WwqVwhI89QvBCZqVaUbJdTAoK/D2Z/sUFllOojngZNkVbsF/69CSGaoULS7
8K0pP8vZqTXB/T27LdzHD+sIUsKCcAp4PsR/Qu6GUYYn7zeEOFMv83hyXCz1dyHqNY/bU3yzZ8p1
KB+RbctxKtTj3vbMpQy1egBXmqIbieowyJEBQ3jeMFNfFYX1o9h3z9Ry31mhfQphVbI1BrZsbFIV
XBKyiRqa6xAr6eDXV2dxmqjqPswVVfC6H3Nqt904H3h2ajjeCYwkAGN5LlUNh1CBRFhv1goqvW94
Uguun/IxphDgOcoNR9joEgizIYK//Jbv4u7RNCg2YeUfP5nzAGP2fsi2g6MyYDObfElOY+FT1qgK
Eeed0hZ+s1CqHQp2WzJ6hqvtuF4v4r9DJOlb1EKeCVpc10JefJNAT2XgcnTtz0urVQvpIivuPME0
kQj8/wyvJpGpb5OMnVLSNnObZaH2hoKdY9asdS8yGWaXSD1kXNB4aWE97V6SRRi0YBAaPJNRd+vd
BSiiTdvyaCNQwapUtXuAF/C47YJbpSIg5wPkDleSE2pinQx3vR9o4v+1r38qQo6+D6wIOdBPZnt0
KOGs68tcFg7jEbXZfNN0FQFShvgFYlS/mBM7bmGO+Au15NmC6FymMJa+kdrwmulcnbckJRpk1d7r
Crz/z2ZX2XnBGJ1F0Qm/uIk2CfKkyZpFK6+7ysllewLlTLoir17OHUd9muZ3ZZeeFxmphm7I/ELr
vWVp3k0OAtYZy9XCs3Ct6cgjjPOLiVRvKb8uxcZzyJq8Yi/FS3h83rHoIUeGfsMKGPdKjukUS1hq
/wM/VuHzbtcOZBgbj5Y+Y7X/GZQ3pZtS+ZJv8rVCkDZinJzS/5X1xV58hkiEfTpkSI6a8wWQAbvL
LpiJwIslG/7fV3fGylgX1Obczwzaj09SszuCxn8BRewnyhJad3ez5SSJQAHMiunAgoiTAkBM5SD+
TLlAdSKdILlOTsB6CzG3UQStAcixUQII9kHoN8bdBz6LtIcVcp+cXL2FtTLLSFS+gsotsNBc0PPi
uqKEHq/Lbj+NUZ4FAOoUwiciSnOo3nQPKqD0UKiMvauAbEa2l7E3HjhTL8NNgOY1ssF1jni9PGt0
qU6EXwF8iHphzjhB+rmZUY7koGHKEU3OEM6wYnMVAo28CRqvOk/efdhkwv19McV5YvA3JStkeNjQ
w3fZrYh4IZ0kBfuNp/mFViSKswpebF/VwuJc9V2NzNWeX48uZuqg1IKgPAwM0QQCa12jYMhs01l4
yeZ+yj1hshGBY+IomBZHI8iissa7viYQ0pXQ2bmZL0xMG/IxNpS4jDG5JlU6X1lSo8aQlkYALlEi
uDDgV3MI0/Ti5dGEEKHBQfyDBlDVt5eRPvm17adsPAwOr+4nY1cD7K74t+9rCXJYPfVPFKJaS7O9
2PSDR98RStnhCpEOl33bKAbUIekSEWwJzRr5VbXb8t4t+M0Bk8S6s2YZrZQHW2TNfmb/VR+5H0UP
I9VVIE/OgYgQnUz1/RWinnharrlNxN/lTM6rORVqA+rrSQIlg7A70jXJP5tbTlTm+DvgRmJpKKcP
6otcDa1GHEgYDORtK5WgUGFA8S2e7umKxPA1hGcnRy/Zks+Z9w7V9FxgB1CwR6DGHEFb3F4IMYA6
7mo2kpPj82uRiW5NZ/nFbzSLeREbUTf/S4iZvwT/S3f+c3zMdyVZKLavw5lN/zLVsz6KxSFy6HSS
vq0U6EgtwHXBhZ1FmaEXgVCEV2q0JWydU1jEYrhJ1RkLVPZRDT6b3aG67HhlfzBapGxn37hRrZhE
F3hQTFfj0Np7jnlueG3YDX90w79hgDp2Of9E8fjoYE4a/o+M6X7ZKPD7DREE/te169jqMuqSG0GC
wK8BeCf2XY0aM6T1+mJ+4Jc+HHdAxi0ILn9YwrE/QFjn3g1xZqSyVStMssBe3INmP2oD/tn+FgW/
t4OtZlz9mP6MBL7BTp2T86lD+FbbU8+GNyWjUFhgQZlzipqfZcDIA1qFO14g2IyNe6RxmAUxRDPi
Da62DPGgCcgabTklfsfsoegh7ZSucUdHVVsgrvJu8tsRlO6zzrird6B0/fTDdRejodL/I/KL7Pnf
m3XCWfDg8al3rpHQEbLjDt5L3wBns4vkDdLoZuvHYf7gSt4tWnz9w0H8IC+GPe+XoN9CPufj0cIm
jXXXsL2e8MF32xGpiV/EVnW7or/Coi4keTlEnsXHSOua9vlxNjqQec5IFYDldtwFkGHcyXwGtOar
In0G/GGH/I3t0baHIiFRM2xhrVgXTUMj4j563O4MYui/+mZ+ZUxfJ/CkHJIlCpAT7FRoBneuXo3K
1Ou2ukg5GWw1Ut3DHJaTxLVfIqtcjuq185zyO6boEhablQ6mwgm06fSCLijTwIPLsB1DvTp++N0Q
NtAxl8AHvj441eCXK/YAJ3MgNszVIEUTJLI/s2BAQPRzHOAAx105dAeOHvJj5ET7nFqHsrd9hXU3
dw+Xwo0ZCdD2IUT8VuIvPd2dPsEw10XuZ6QadA0b8vd1H91vSCDlzttYMQJ3V6jmjCu4alNFX7MG
asJfjyHlf726qCj7qyNHt3MRYZehqaiAKtOoJX9qLzSvwFIUS8vzMNCKr45oeoJXpefHBJgEtbyd
RRlGPa3ovDuEUnarHLQpDrDW/yU1F2WRi2ReWaeYwyL8piW9zM/SQfyflIfiy5FQnI/HEGRZyi9o
rQkEMM6o7L/XIrlIgOKQXdYpcswEsQzs0eKf23jWiEU8bCrCiaxgc3MX38lvKNncaH3IGv613UGb
fLb+TTB4zPkdWIHA3mjcIbkXvkL6Cgzo/QUx3qePs8aYg2ozFj6kkaDXJEZ5sOO7sW9eblsU0OH8
zHiemjt0YhJGjrhPwjmNCnX4dv6EcPY/aPvF3Jn1gkIARf/qspx1/ZKP99EumMHjt43dZqIlKv4q
kZg/jDz9UatSF9BV2nFSuZH6hADJg2DQCxH2ME/M7bxlJDB3c7PIfJeXl64//XCgKkDh5R/BWGup
IHH220yTSMHNcy3cQSF68r1a6I7zu8sZ93V3gD4GBi6nB/NoRCiAsJrZTWARXTgqWW/bKWQ1zrcj
152i+krd7y1uH5edeMX2ynQrS9IrXSU83T0y2kn7KFf/U/0f6Ejfa9GKoAh6Ua3GKLHHu3grb/CN
C7uQEOuusUEKKB/vksDTn1N2SIOsywafOTYQ+TcXWNlY3HIj5T0T5RSgDsHQYa3J2TvOeO0zfGLO
uvm5U7dRJQ/r7YcNQ0mxj2QHaGu1nQGPpBdVA8TyXDONi3VK1MMFlrjQCSbPM+rx2/L+q1jBRTfz
vRa/vEBVjJGVh5vGIHqr8EQh7fpb6pYX+UCsX2TF31qy9TI8xOZKHODCgJFrqWOF2jXUftT8rHRJ
fjcWEBWCddzxGEKq/xVpoQ66PBMPhX2knc+3JWn/LfAd7sRN/2yNljZiHX0A5FwfzkQQSL+OjTLp
EKpW6kOTNQLgz30qFwJ7QCzqkEJgYR/nrRfyrHjDEDyOA3cLs6lfn2ekIYAOnQCBAKcceb0jLFc7
O9LgBPc027+32OWxHFzXtz+mZ7SZJ4mcV1zSQ2XLtF0wBSI5HR1HVkgW4XXiRRvTKvwEvv1Jr1ZD
cm02OpRJqc0WTf29FTKqIKHr/DEC0zjOAsrYfhkrgLLWXsSOupnDijvmZVBHfy5uymwPVrT86QHV
KyUEG9KdOz5KdZtjXKGqPF/W3sIlALa6WB6KT3Ma4JMjE6rnMVHc+9x7obStLGdDS0Dt0MC60MhX
g3VVkjt1y/UE2GZJaAUlnLH+NsW5295g5OlsT7RR6cdTGkKbJ+QsjxE0yqWyZSq09Yak/SrIAP3E
lcRdcg7ZK+R86A/65qAopxqrmaNTU05Kb5tZt2eeDS9P7NCaLYH4k1zkjCkgfPWPt0iPu9MpUsQa
Sm2a1aYHPEiHg52BNzdZ/OWr7VDE50Fw9U9s914uYxFRqhVWoP45r3iy0JndcDSsD2YlbjyqSvcg
7SfS6w2ty+BXBPBv23YmbNd2q/Z6hQsN5Wl3Aet8e72F7Z1/LHi/2kizUIynZcdjIk7RY7TmTqxb
ETV4cTodyPFGqlIVMgonahYaxxs8ovrrpzfjtdGuTPdgb0o6IEbyFcF+ZEtVH6tY/c9Gl3Oo4X42
1eEsBqgZZt3Vc+5IICYAh9G7cd9WSheFMp44QNnOfRkBJv9OJnka57+uG3QWacEr+K52uIo86jTA
1M3QiL9+ZEgR2/+DVZPjVc5m2GrkXmZFGj0KnPpu0uTWWblev2rxkkRioLBMwLKmbzj46aI3THG8
2XjyzCqdBa/+as9Yh7eOaV0whfxBT5bLIkrPZ5cZBWj7suK+6iS0hnWHt9/QIIqvo3RhAT1Xsnf7
/chNoQvCotWg1QyO36EiuHoCW4ex9v5UpmM1Dn/EDxf2yPC5sq5UYjrWmwqn3QK5XDCKJxw/1fwP
lMS42ny1rjSuMU5L4G/DNrWkJHdFrAL/yrC/wghkQkxj/58Tc2cRs50xmaOZJRBGBZ923CLLd/QY
eUwZS95PrLI0GRdZlCzN+qYwK57WBsVsD13/J6bpuzv+HMUgJPfblbioCM4XIpC0IiVssu3DTS1N
l5j0MdMKxdDgaIQXp+5sQmKx4Wgr+zDGpfjV8l+oD0Z8NgL15RR9RrUnNQW9L2qv8c6U1ihsg0q8
VL3v352oM6XZft0Ra1my8tT1gf7hhgzdJt/gzBdUJfZUQJkxOS1EJZbXXqOj3GCbYsP9gZ9Jgq9d
cSsEWQf1yNU6+72owgvTBjIr4mcU/BkqPPXKYeBCqESPxvBR5mBNqHdj5zNbzmLgauzQYWiLTEbN
nBrokg46tKEhV8Iom4sJBjp0AeHWSOjs1NHhZZhy8CTnYGXxe6N3t6rPRGYfbIMm7rB+996AmBds
MV9tZKit6NTqip43ZEPnzTDNFpdbfDXLCv/em+gPInHaD26nQYfAz2KenRkQan2JQgktjWBMJL8F
9IYNP1iM99R3wbCkxMiHDvwAJj2go2VwiR+qFNI+VicLauw1PJn56Fazk1CGgu6FmFuAMzKMEx64
RhJmX3J/97jn5WouvuIkS/WP91nCwj6b5AR5jsuiv7bAu4I+PyPm2CmNaVU+AauPkYWqyqWRhpAE
xiVnhZAOD4IZP4O/7iNsGDDyB+z8RLDXs/k2RZpkRit/xGQd5Eg5x5/rNU3IRTKcgXX9fMZuntdX
XwdBIaR7Ydpuzwp4XxzDbU9tZmwfzix+k+BO5XCqklqL8kIuSF84ayBngBpowi4W52rJHxovTJHV
PSxv0I+0lKFbVt52pf7gP1nPpXP2TILf2Y+3o0qUa/eScjK3Sd4T+3+K3a6PPwfrQOkfn8Jz6Z92
ijoykVBp6fodgDFQDxkMR0WBTFNwyHlSiGR1wsZbZuDsUgj1Yrqv+QcKiZbWAj80BTDjGSZMFEPZ
z4HBauzcuTADv51uPP+8rljgkt3D22O5WcjOPSrTXXCZtTo0u2leFg6laMK4GsChZ3GMpaMOaifA
3HyiEz50dYYzBilfDOGuSEn3ncrs0RMaXqnC+1ntEGKFG981ACJPdAh4yB3mwrGTq1DDd1AyhymI
WdbRhs6F+kyEx7hr4XqFTDW2aJgfSOMVWk6ZIUKugSd8MmilMGL/ieaWBDowVclljX8t8h7AVaVN
NAdPqYZ+bLk6SZ1KT7PObdz3zcBgm4mTyKgjixCqeVZ7azxObDiSF/YOHoJMtQdGlvPmVkW/U0rS
no7gJM3kDwfkEcOCenStrRiaSIFLxzySvhVhwipM3IwvJAwbo/nMP/9ktNUvYNF/fRJlhs/uYtGq
IfPVDJ1FFRADEinKMe7G2cXoU0nFSaonZmm4alwoDRTEn96k30hxKKP5bEOEcZpthuNHBloAA90a
lY3NJzEVEJmizaN7Lp/IJpW1HjBMDeXK/Qun+90kDWwLVXl2J8XpPIC2It/pYLE/zTWd9hEeydj+
bkz8qxnn+uAG1WSJFhPrZDYLKzXgkQl8jk9sxmSc++1r7TsPQtzghJo31BAjYRWSf3f9nwbxtX3t
H4KTsxjcm+NYanJceheju7vu2Zm8lV6eXrm5d4RHl2Vhx6nlJdUX70ulYmjn/+k1V8ZOHuiIfudw
rLsw3G9rY3yX+FIXqNF/AGD3+Kw92N5UY7sWOvI7VXvwSndV2fw6KzoRUALDO/I3Ch6sr2E5Cvqf
LoGHHKK74Lsp7E99KonG7oZXHfsw1oBceMiuATfeWK4A/wCBYOBotTJePlTl7p9saRjDdTjBzhbs
JRcU4JQ1oD4jC4NwcBPtxnNrqvqBKrTDhOqF5UTbzPkY5k4VsmKv4QcMjFBsf6DOSDLfNtevC8z9
hTsZ6wbn19PnW+u4xRBAbjW+wF4CZ0wZ1cpMLb1koxlCfyDRuudPjgPQKiiQesoS7TOAFXuEMrFn
3uFriTfKjZkqpNPEo0O3EfOfHvldstIARlRGN8NNdt4/eMtvntoFtMI6FH1HI7CKXCEoLdWfgiG9
OxyrHOzVGhRuZ5K/RFiZvwuW1HDtLDBce+CK41U4wopWzskKETXj5Vow9cUJ8bKhYoMINSlD0OcD
f3hn3VObYJzz2e9U2E/dtR0D9SdVboWM3fglal9U+dYXLmZ8+3wRj7Y0LWw+Acr9aIWFMt8IXrwQ
eMNzCSUU3MPrfx8ZaM2lhd8O7noKSnCDVEUwPXs0BRpKwm5+V4CVE3yPSMVge06Pbv155NWrZT+Y
FrgzbLfW/aMTcqfDqzDfj+0AdlEVnVBAja2lTKEz+oU/42GtYPKvR/6W6X+UDwxm1zoP01Dn7Hh0
nVN7e5YRHcMiDnwacrB0zuNF1pshW1m0Zu4KN9u1rERQ16vLx2DdtYxQsYvrtL1lN87x3dMKROLf
h8gWc7o8uofXLrYlTKfnhNNAVAMkwCDe9DeIqm9XQuI48U0qNkvJ66SqH1CE8gPYuEbLQq9ne9vX
EF7RE0n++v+GUpErB1Nz1f4DqBHkrvH/Y3Vw6Bh9t5ZtcgAxSdUyEBguY5Q5I5DJQi5A+VB+ik/3
TQnY7HrovQJ/PlCSsnPz3LWpwrAgMk4KaWdBK1yIKSperUW20jlt3dlErlqS4d5cj2nG8D9f6nfa
KHUYYU50lpKGVjNWLLhwFIPa9Pm29Uu0nF9V2ueRGyXNyP3HMYak1iXgvMqmkBAyrWV4keGF+zaR
N7EwZiNIzT8JwnSk0g+3UwEC+XgLBBL7Ylf0S4c9hW/B4vRFNd8JPK5S5guJXYw6RK5uzQl7iMp8
yb9xAo5Hxse+/n0wOwtXsK5NZCmb64/5q6JssPCveRMBpCMXdTT0/06h7wlTcPoT1wrJTm8aHOSq
EExl4sD4RFMwjdbTsPDqcYq8DAsYzd05j4n+XKl9E2MEjwRR4bFYEl2KzXnXc8o+qoaG8tGQE/pa
HXZNUH7ZaMJZNcDzY/Iotnsl83OdsYQ42LpjDkB/6sh9ElD97NCOwe+FDtc8pyXZJLeoR2q2lElY
nfKkewkSJ40h2QL0NFmaggmzDrpUN9lwqZZRNIBjJ5zKp6lvOkK3Pj9W+0KrDjMVMiYfrJGeDg/Z
SBPznnIjNkYkD1tziZ4kRD0gFQuszbr16RGk194vK0cpFklZRWMWX+TqPkhMmY27Ur5Ueb3Z9mlv
rmxQF3xoydKW5eGUflF9woKEymk7rg6VKdoXQJglUTDc3Lf9lpVfwowBiA6O2MucCEYhdujiIu1e
bKogI4H95dTOL5U1dTazyJkGs6rgZIYSwR+E0zg/hUf4o1hehxBk+RL1LjKuBK+go0+gmjbKw7m7
KcncxMNpSFfNVdETxHRTlQfyXgadSmSFHUisrroOV43rJzmo7rp7TPecd6urliMlLltTr60a0rHA
Z6FBubbJXcs3Yep44HWFgk++ZgBBIxqf6aIjUhWXZrDVn/B62af51jT5mZkzQkgt4vftkOH78AtL
4zxuyqtJb07qjRlqRhJtbwJnd/oU3Y0Ro68pAjpTwQu1v4HvevZzH7IanWYmrdX+ZRIsYPSRdE84
pLq2+CFwYk5CvCmq0Z/BcwJwwewjbRms+Gwfo/ub6kaUWcOVNsiYW7Jz6u/8pabZgXGRgE1kl7eC
+EIaFkVQSaCA7vI05A8PXtPt+cND9Th72rrubaBsLSOVQKn7++SmxSJCyXvQL2E6qHt7/BnH4ZB7
t7zfbfdolHdAPesvXeFETv57dEhKY2I9+goR1tX3BPM6yn/JEXIlHZI6zzaPx+ZU9n4Cp7xO0sYC
0vtHXTpl8EKqTk6RD/3tm9JopapLDgiKXALVsIFrfYn/Fqzf+eQ4kewqv2cCLopkp2AFBATT/OBa
Ge1V1TXw06AEvFQQmA2aOlpSUt00OKVE+38rPYb5p9RTKcJ3E7KIXmbu/hiLfyZHqEjMjqBUpB0f
0NFzABUnhcW1c2/W0DWqoXGywUFehowlL01Hy2TEUAIChnJHj2+ZPzMi1njRFgFtrbo59ewC+Yga
nfW5zBNY2j1wuN0DH/YHEjMl4vlMn95WD2X1xyNXEKpocDm/Hmg467fI7jMaMDPzvOPjRCHzYUtD
TetyprgLKMiKUU/4HeIrSqqQVfiRFY+CeZM2mDUZ8mbsDr5Z9O8c+q46m0AhGyeYy+9e6YwYRm/x
l+kd0roBWlMQxrVQStWl7e5ZrM8h52kRp0msgJ2kLzH8iK078emuiNs/A3UAq2Fq/a1GhNCtIix8
JdxeH4+qV0jlX0ygZYmA21lw+afhc36hwHB+I2wzDWTcIQXmoN6D79UasVzAE89a8Ni6/L/asJnG
nvE5L0seMA24dgFmDXyhbQyQh4ea+T8LMQwobHLyVdIgwjQK4TB+ERSIDoT/t/umnz6wivQbRaT+
qOMdqIbscvgfVJEpRTphOzvxCVUhipAfLHeyjSuIJXUPLnEnZemtNIPelXQRQZSLDLlxBSGxp0Mh
kK/8oujJGSNQ98KbXZKGgpU2b7Xg2kP0ZEA0uX14dBvJ1pOIoC2zxQaFp+UDAt4qePbHgr7m6g01
j/nY9s7ITdnQSndO55xGgIWMxky7HmUSZz0hZBMFVkx5saa1dnurSxT5XV14pZTkxzVl/n0HTaxr
6fiEc32o4plb8a95AiXvQkzUnqMvdq5Gfj+gTckoHwHwrbJDdzd+OmyaLYZ+faAjHZatYFfqgsUi
rKyh8F/grfsrFqUR5d4V/kBvaZac9xFHDShIs45FFKjyCsSQC+B9Ipu8G3LUsyfgkc5vcvHzlTe9
tVNA/VjQiCstNDvXcJFLWsP+ir+f2wsxuVuywrV9Nrd4ZyaWXfr19r98tm1uhwzphHUYj5OPIhjE
GuSqbZEPZ9RDCjkgF71hGurrTs+//qkDNMpY50pPtBrcNqxzM5ZtzZQOlm5LpxP2AW8oaFR757Ag
0O/mc0f0KfTZtL1gsRPW5dpGW2JweDw59P91Tbcs4+HQhuRoQwfJ6qcFupsDUx16iuw7bL6sqXOl
IXQY1e3j6HgmQ7B5Tyv/mpGGvSAMBjQ8MD3uwvOXd/tV0OC+ArVtGsgqdZfN/aemslyrQQQHlPnb
DjpvZ/0lsSZdxRwDshM2jznSUsMEbYEXsascRV3F+WhJmbvrJOPaBQcGuBvDk9rAjno2blg1QNuu
NvSAd1ZP2F+HahO4V32XBmuqS9nt35UeWgF4fFVJLmmiNtTJM4Ui3Plb7+Umtm4nAJvWto6S0b41
eJLwmwedMvBdUZz4uqgOfShxj+ZZ7ZKrb+4SYv92dEWFK46jLFVgi7+OCU/RBFG/qTFh9fTdwg8m
s6R5G/X31MPySkoatKQMaKDZsmb1/e6DwJqyVgfdd8rJyZBOcjgINQYGZkt1bmWqyjS3uI+PGeX9
iYDNUwQfhEEogJBYhr3yXRJwCiocXV32KiKMfU6nSQl1CGJUHn7y6uZgrpZ4Fa6TAZPMrPKk+088
5pVQ2MRxUVxaDnRwOxVwG5wkfF0k7RwN/FWTjiM27fV8rUBnSZM0crLWsX2+x7JPxqoZrzB2L4Cv
001o78py4i+q5BaMo/HppCtu95rpExGD15RzJ1TvhC4hmDSLKSWnS4+555vDojDdcqWxg/plX71e
fB0niTGOiDC7E1haDcRWoBq2wuYdvhv3MqycykepMUVmjnIizsv7EmYJHpnDC8GjaZwJ2sx5b/fd
aX3oNJfd97LvlRYOznfCxPW2+4wQmG3djbTNC4pBXzk0OtSz2jQdcfN5WQdGg2Wj4jRQ46UsMsxM
oBtrQOpyIjkM+q9R6a/ml8reqto9R0GXIaoom+79YBoq8kbkZeCZ9mRCzizwvgPdqm8GvXY50aZ5
lODCctrri035IkZ/eKTYY+rrURit5bjaWTDSv7/pav95rnchofR0hWjxVL6jtnKKmnlgax4Bmw1S
mbZj9fNp9dG9xU5rXtdlbNPpF+sUdwonbzbTonzj1RNr8kFRWukkwgEHYvokGwQqbTSzMVYK5vAj
jlirziNz2Hh+IiYjjrVHhrpbs3oz+kZsghOnW4HmooOXrbePst95SnYadOZrE+3V3uc5Nzm5TMZD
MVtlV1qt3G1NkGLHjXMg7GSKDHuBkS7X6M41riQ89+wFVEDRJFryzI3Gp/QsXAFPx01YDUp7PIOZ
L7cZF2LYYPVmSyNTBmobbKubj1lLt67vSJSPHADF3M8129n7ElivyGOxeCaYXH2bYMCzQFa3vbnj
7ZVKT5/W5go1dQQr/1Gc2QIr/IvxCyEiNjIweshgXZLt2rvVUXtsJhzktndH/oUEtAyqBqkbjj2J
x3OyMqbsz6sRcQ25GWQEg6xOgzTF4eJljfcVzp2lCL2QfKyY8ZA4NCY5x/7w+nH6YDRCOuM1On9C
PxUBPJ42W6Dc8lxgegnvBOvQ7afm5liekFLHxOIYdo5cOKdfQNnLDNvNSNsW7/BluCm5NPrefijS
8DzJvlg/ZBsmgbuKxdt8o5NNBZoBkdRL5fzNgnOUHENc6m/7K6jvCcOe6R5e1U7+uaAM8HNRI6Sc
1N6kikM1bzLPovOSg/lvQB2Dls+FXrNmnDQ8Ls4GKim/PyPzsCizDtUVGSuqe/mMU6a/YFsYU8o2
RyX6Sc90Q+SoMGNG9F/hDe+RpfrQOszKleUHKw8UgDVT0QwEmRiJOCMK1sBbClJLQaFKjooR7kgv
QEwf9MD1/IrnCuFm4Hxw1vGku/dMHGk4DDmUGdjtrEr9vAQhLsksauIppzac0WL+24hNJ0NFkQ3X
hDAyyJvo2HmrzsHRwbE/AMCUGrxHrXWBUnt4quPPu6+tO1gI3+lkfSCFJWRXWaZi6+CuLW6TYuC9
atd/jWHR0KkKKif5GxAK/L6eaKcqbGrRHFoOYJ+U+0kxMSkhf4Yapl0vReQJOh7gaBITTjHDz2/x
nXBXlHuiGMhCanCTh5SuyjN2LwNmntjSh9HBgczgtq7L2kxe+vlBgywcYAJhXJEUp9MIM1R6UxhN
ZNjq1oh9C4Fju6muQHir9BYxvc4loeQlC3e+iU4EtPW21UQXCqVNIynJ0CKMyl9FhEbVTkOvMK1e
jnHVz45xuCQSRloaMfQj9KwMM3w9OKrgoxO0UssPUFIB8V1ZcvD1yjAtZERcJ27NGtdK+1OIXN4U
RJhk4c9LuIXT/FPeY509L49KK3fW1kPyOsdvl0bP0FoDzRXol5I6tUFSA5fVih37V8UaM3goMvO1
fzSnCo2EVjWi3R4vAbWNB88I1JtgoOylZ5M0ZcHgETGYat5iuph1q22RxvVDu4LgXWLKdaC3LrpA
MWIYGaKTafecMHK0BdOvPa7L2iY6m2FMPBYvkFdISIhlDP8lRK37kbyutdWCR9K1PZLbOpsARVw4
+1j1BdAozjzmn/qlz4H/YZTLXZEoHVd3eP3Msn0bDy1VJrQSz+EgBU/X6GO5bPd+/U/YF5z4ybV5
xuoFgPdr7cA6u9gH7vlldIZ+NcIzCkAb6s/3ecOPIKnl75yoH6Y5cK3bOuD6b2BSg46iN6dlzIOC
uHuTDlsCr8Bb47lTnPXugvenQYpX4b+iVYlNQ6KdmreKmeyletzv7ZqYfRu0jkbjf+XQgsm/DBoU
X8HHsAv3ErGyR0smofLwZx43R9kQhizkf3Y5MC8W750mUBzdv7O0GdMHRrv8ua/1au0FgNfZIqkg
1ITdzMNiQ3jrLSHxQ6eY9uxiMtsYuYDMSDHdKkLa3pJKVxLYE96Hzxi8Fj8m6IZAvcMhrcu5/sOc
Y8tu8BEKFsv0Q9IYnyMo5SBbOG5kfKeBpClQwO2ZnI3KKnY2lUoeEzEcQ2pGW96JxNNybhyLjNnz
bl2ZqoYJ36yGuIEg84fvGwzxlAL6hgz4WOx30xvmLeijr0LwPoVQfncuhEYAsZjSfw+poh9j7iLj
nqQ9YXLWkPcvt7hLu50sgc5ODLXfSjfz4GV7fSHyJoft/4ne/TqWSNAgr8gUrJnTDjlUqADZUpuX
pFlRegYpAbApwNSAVhN8Pn4b7XjWuapUiod0O1y0y0li27D9uNrxhriZLhISF2x8qmVgPL66oXcc
qf73+4woVZKicYIX0IBwywVJW+0WLLxJ3lNIoSO6NGyb14QeerP++LoXFdJ3d9n404aX7f0BWXBw
aZ2kv6r//MMwaATAK0KOdMcEnMAUdW+8aO/afL8GlZRi/hK0eexc3krP0sN9bUOb3bITrFWv/2Wn
ddsSWBf2bR9A2PfLKmre5TPPsZ7G1/YonSSrkxCsE1R2yCdcIVp7Y3OgawfxJ0WIK1iLeeGwnnl9
OHCk5ItdXB2evF4LDoM18gCf5DEMFIEBsirO5BWolam7S1MLsNhojKkaHbvaSLhaLf/2E4170F38
SMY2MStigxKzytsUasi4RpTMy5qNFbRMu5nmm2ZAeGnmx4hGD2dPh8Gpf6PebeuDWlJmRAycH/rk
U3NjS32zVGd5GaH5lW2sOKbsCSc1XIf358jI+dHLSMbw7IqEoPJ0qbTJPQfQSC5BXs8uacLogAkZ
ezSVjj7D/grKqMHsydQ2jwMYTYPeaGRAdDLuOUDNLIj0O4oTyVDH6KH1s+1Ok3ePqRHzc7BHCUEx
6eG6Q5x/vZg9dM8n0vkBe8B6qLHjrHCUMiySANoNT105B21t0kaszePNBzePP1CSfJM7+2pLLmwi
liqIHd3xqiCGuaxDQMWqgM/iNTCUFR3XEGFemb4vhJzwC8rZOW6UP8uhLlpEB1spI86zsz0v6fqd
2jno7IqgjRp473fwQwU9o8nwjdN/SdjwdQkGgCYmLe+t78/YB00gpqNLw4valmoqejP48xhFA614
WctfibZ9OtRpwkVeLk4tZHHYjRN/u03avDw8svCrn45b5LAcsl7Gq8X5W8mCuwDCE1Uoov86KHIK
yrl23JbPKD9WFq5BJo8UYOYvKBTSG+twQZ2iHNr1N9IkdLIWc65nf/o0cq+JoXHRAXwdIZjQisi+
Hk/Z0EyobPWJ+kpzJd952HAsscMx0IYD6qI1UA3zy33JFe52Q+E5yytVwTtD+4u3D8B7SlyMj29B
KdKDbh0BtJ3qaIAzfFzRF3Rpd7E/48OWMGuK0myOppdXNkyksGRsmBDxWdCshbtR9X+YzSdalxwp
uVzbvQTLtCQ/PR3cUcNmY/87O6D5jJVwkhV0iZ9r4UhGZ+YKsSrLWyW3fmt+ci0k57Y/gGV3LMgR
OQmfIWvIsUxHopIqwsem2vyuNCFcpaygXeztx20dy0cZYc11OY24KcKgoTYQpjuSFcXxb/VM72Q4
eUd5bQRrDyRTr4xkssIDmQ0YR07guqdaUwfH9D6Dk/n96oMyVGuDDZTOxDHTeBSmbZOZINphiQR2
Mc99d+tw0H2Nq+SzN0lBxP8b6CeTjrEoRi5FrvaMUsbaGTZkirAbD8KhE0DpWFu5quQhtP7AHdQ8
i19ITZQH5DbKOgXPui8tcJ+Nckat/dVtCYfhEe3V7r7Xclh9UPn4hBxa/+oImoXLwXtUkrd6b1w5
dnw1mu7zLlc1YtK3EPzD4jc5q5hrUfFMu7OGE0ZB9EIOM6SjUtCJS9vL/C3Z+8sFSwfiEnNM/uiq
1OzPHZSj4cJVd68+vJ1ZVkIYhNUqspGBQ2GVeYyTTdJP7dsyZEZPdXGPY/5aeUmw0tUbMOW2l+L7
2aMuUM2DtUGT5155YPjH+GLrOVi0TidSuUlf+UhiKbNc9r6KYxMRgCgs0IoTYHkhe8PDgLpos40Z
lORfRP7VbAL2BFMleqNOHBUc9FUPKLMuz1viO+s42LPWNH3nKeCbZF8RsQADeskBTRqGi+3hldaK
+szwqPLsHcTwEc240Kli6slU0P7TIteQglEcitpUIR30uO15ZbRVz8nTpQgkVMba8/SNWpC/+cjS
6VHgHDj9Vi0x4Gi2pOiWSyWM8lMwFxa4ehR0ZudqlonCfCvzbhoCxlV6soLrtydGhVrSC2L63aRj
ulLNxYj5wqAakwEtzTVoiEJJVxioBure/5x4R1wQJs9jxPWGvF+kmgDEPrmqZEmzd/C61Wupy3zr
zEpDoClpxAY6Y9r7BNraVJxKs+bkPh286Jhpz7FRykW05uqfDJGvzwI/C4JomeMMkumXzejnDLQD
5bowgAUGTNofwzwwI9CCu/EwnF80/T2TN7Td7wNITS6/9n1UcmGk1vqidJM3uIXMjN3AZkbgPaR7
XQRlQP+bTTW3PX3U2Pm7vguifquu3N3EpAcm8CItjFgEPlUoAiaLfXWbbbdmJ/Uf7PK6s8Ld9HUd
Z9SRujtkH1daHLJHE8dNxYroQ3Jf6c+6KmHPggJ1L5gDxeTb0nfJOHI2oB+N3MPZmbBkBhSAitN1
aP3usfan7UPtOWy0ZgjwTPbVfwdJvYMSAiS8EkTLtEaiAvP56KKrCxM55IJ4ITT1T6Y8QPi22Jrr
yf9sZ58Fmsm21qwxhxQQrOnZs8vUlnWpFswWl2kUdrX6bRXQuWDO8Q86GF1ZMcme+q8Rva9nPF1m
7I3we72CZePCVdppH68I+FujfK5pTHoZUSiB2i5ZnVKcKRRgeJmGZ/swgatUBCz3MRHNGJdBnG6v
0WbDsH/G0yR0e+O2oE6ta8R1ryNXXHy23bV7jJpQojuWDNqKOQopTSEL9TlKWEX4eo0G1bTNBkpx
GuUcTu34btCPXcJZ7hrTLoAL3BWNgaV9c9ls6WJYTQdFyQCIXaxPax3uU6sQbodAhNg0oMpWMO0m
R3P8yg80CkRA1zzUu4St1LEyw/wYvK4hrEarkLc3pqRnWi2WmH2VbXtABJUwr2BkvQ2YrdTpG0eE
YkbbWlbb/Wdn4rEFApl3dBMM2MG8qEDUfsdHYhuSplUDYtJ9Rn3ULcN4KlNxtHify+CtkMFG8oLX
+jDDBBYpAerABA0yBRtUeYI3Qd5MgiJanFqijUiYRa93FomwZDMBy8CgFbkoWvLUANCN6P/Of2+W
4Z8nM9Mifnu2AxkCF7kuoeF42/wVITMAztJ2XIbS8F3f4lx35Z5E9E47b4e912EUxEq3v6JG1eBf
dY+mMzX77OQQ1Xyb5I/cR966QgQqq4LK9irRdGiouWuFW1ma/a3ds+LWASJnJXJtb+V6n+9B1T3e
wRbFg4gv1QRSKY8GRSB1vVaWtuP2vZQkeCKkF39wVpEyJUapilw5sVkiRVFOe3i5FEbztJxKnySs
hK9yfRTgDwPyOmEJCt3ZW0OG+YvSGKQfVP9i0kk4KwRav05p+NPOAyfgAGzRgeS38M+SPaEcghNw
e0zL4A5WW/kgffBVqI2aWURxTjCthMo+P+vCowmG0shYMLXrJAeufYCyl82cFqoKDNv4Ki3dn9ha
F/WctsfGz9S3tCLwtEAqL/L3K+PKTUA4u8zmzHp9keR+ck70SRx3+Z5YidEzTalcgwpNq0i98l2d
KfDi1Ad4+NnPSxLDCw/y7fAG8WddQrFvEVGojSYvDbcZ0E6gKDqNfhyI4zOq88OkyWoOYHvfXu7C
IPkeL/xEIRDfIUnMyRaO21YgSWc65q4f09PyT9siB/YbptDO+DTerGX3vWx1pied62JUjl0ykM7B
KFMQxQ04UAyQ4zmqIgDfeogFc7FXNWzpD48XgMOYgV7iWp/qJBggG+LlXXuOSGUy4GiHyxMFHFYT
Yvn8S7EeDDkkjlhzyAOoHG/QmIMF02Rb9q98HX/3UeeL4MMKKYUAYyOO22TJyKA3dhk3rE3aQgS3
NY1+nQCiNnIEt1kAreb1ZWVV9io04+EqrHWb9McRzvnpmBflccoILyjpLlCCZJOHnjUrN9L4Cx1+
EbrbGG6URambxwV7DEhACoLB6MmxLL/lVfth2PBbJxQ8ZA23jHHVG/wXXkYaTjJfcsg3xnJeTBKt
5PUMn8UQmBoD++ObpliygOubVIfmMFh0WAOvZnXzyqGY+IMJ7AoLo6uRSmli7Vezo7S6u2Ej2FqV
iHunz9l5EvOLyKAY2w4S8taO6Om71LVL/zLu0M8zplN4t2ABMynteJAZASpMQMdCuLIb9fmqoEh5
hd01zkaxQe4ruLE8P0FAG9iXo2iNHXCJGUdMXHEhbe0cvMCQjkxgKvkK5W09bJKINlviHNuqsoAw
W1G6EPq6GnVBm8yZYNg7JLirJ6X8OPaJ7CPs92pl7MCYm4QxXki6+/Sc4/9I2651/m22hZkL8D96
jpo+wCF2Mehbi6Y53DtGsxdA7x782LUeu3DYsUrIXe5AeQXOxAliTsCY0bCx2CsnuNUm0G8Sqvve
n+apAuQjzMyvsc7DHCeNpkfUPXNHKeLU13zfQqXASYAmm7pCw/trRpP1QNMqEjecCH+cbdkuV9s5
ECQGTlIs729f96EgUnEwVMONZPPGnsjepqyuIJGeBvAtN9vLYLEqw6GGLXxfrA29sP8qOf6fVcuO
/SYkjmzmVqtUMLFOyTVKNLy/m5d7v6bKPMa5jn5hpLqUtk64I6dvqNZKFJukVAEwLdQet/h09ccz
lMQGBzu9cbjZUJYhxivP6Q3/MO6uAvHBpJ1nD8h/Z0gVwfXi1UIEGccF2j0K8h+G1T98ZE1b9wJf
ql//aQdlJ5s89TEMeEHtxqddxWMViYlQ4fmQU6HyYj7XLil6n99TBuikZk40yqNOJiKsFLKNp7k5
+ocjzrO1K4WpgyqhnA34RHJ7GVDu/ysVOppDUAak9Xn9lhwWn4YmAiau6ljjCekAadlf7jbafy3Z
T2jP/7xmLEV0nm847EbS+YcTadKvLx6UkGvxyP/l89UEPpb5izdzxajuficNJq1EdlbvXzBN4IJi
Dz4r8JA9myx7WkMae0gk2fho9d2JkTAAJmII26adssiMMpcVJLeJAHRwM7FEPuvboCJqwZZkX+np
szE5uagMmKJFT7sxQRDPHzo4UG+0ccGhA+8TH/txYksnFg2cX8AuvtJU6gr4p7ozJDtBYtEMPk+G
KpEJGIR5M2geTmy/Ddt62eiGHqJfG/HV55OCVaeiHJ+gv91+TzpelcyuAoPgjKudX8RxAkf10obn
nXXAbUrY3f+5vz9y67CtBY/t14x2XH4iNSQXGw6gECeBRAATLLXJzOq9dE2VHFikB5KyT/oUBmQk
A/t3cXCfhXkGDqOy+mtIcqS+wNNvUtWVdxrwaz+Z/fHp0gd+PWJEehxPKLYhSxDkBeoBUkMLXbps
j4X1kEhPA7616/j6Lf8qSlhgKQ6t4BZBvcSKLs4xcnMJnH/8rytGvHit/1Bv2/ono8YJwICTvqxm
NzNP1Yz7o8Fxuxkj3ilO2p4XbyjWjGcJqdYAZSCD4DTZRUr1r937I4Kd/BwkobQHEak1PAYYez7j
ww15CM2hpycPg7zDMN5bTPcYL9a0hBfCn2POi6I8UTZErW0cBQMcZZjBinx7clGj+7yjhPMJ4K1k
Emj/S+JlKkmgKskQ163Bdugb+WPz5Ib8jqhOk0xWuFW4AfPwY5gekidiJzzLiOQ/Qrsscx4+fN81
NUUAhyDR82/+5LhmHSsfTlrvC5bOxN7wBoe/fu9ndN9fJrDLGcWAe8oqSpgmS5evKBAcnzNacXcR
Hz60uxZh9NjfIaxDeZ9SM19KH4ZVzYuOzhd3+RRGQsoXdgELWnOJq9JwXK0AHhuj4NprfR4K9gnG
AnjdBmHPvVrwJKMwSj0ihSFQB4C1HwTZcw9X6FAEu5RH1FNGwaYNDRYdlQTSjY+MACI39iI2GR2K
E0A9z2G4pD3YJ/5Ognuz7O+RGEms5GsUZ3+ZUNVmXGVDr5toAFpTuw69Y8Or20B1zpcnxr0uBkjP
8QbO7SG1R96Y93CNw87+QckaYoDXVqNIVxCSeeJVuY4VStS8HUQsxfYdp4yu/pDLbNt9Nu5nDM7g
eixmzA9UcZjqWiIUgI87mjtiKZt1wn4wTrN3ESFm8EbUXGL5bakhkq8JiOEOdPaE/Nt0VynqEBnA
yzVqnN7nTXldLoRhdfycHYzvTCjvviTGv4SjJNRNWv/rzbpLJAUwrS8gJhZI4dXu8Bxn35XTYuqB
2YuPMxPh7Teh5n+4tsP0s4TMt39iXuCh1oRt3N94ZjR8j9SkvUZhkqRCe8Wlja8iCYwLgndASAdA
NjMYNThCTmPKUVWT1Osm9l5mIoFSYmAk6dTf9BOCTEoAZ9Ah9En32mYGScFO8wPqv0DqNDiR9n5P
vbDrp42+xMd0jPeWHV1vW4mUghPckOSmlsCHVAsGa4b1n3fUcWXjZkxxz3IjObTfueJbBYrGJ2xr
ZvoO3S+/RX3a15LkC6NayPj4h54QZ5653aNKcKZPP+XVI80Sc4CYQ5y71VA4YXvmley6GvDdvUL7
QTq7DQ47CU/cqEicdwRI4uqxIGJAlf1fSOa6yT7Is/VJmWiqiB6kKLrKYFcarvBEmT4XxnlFukEg
mlHBQLeKFGcUhErssXB7F8FIN1GV0ZExeTf4y7Yzgdl84ms+giNNaH9iQQvQ0gAd6cBg7jeVY5dq
B8VSc/STe2VPL/rUzsFGyP9DpSNAfShWRL3IR8eJ+4T4bL72fIYYWoQ2a93eQzo2Okz0Vf6MjPAJ
ynZqwYu6KdH8Pv+99dbYPt/qoYB46T2GLTU6GSuFW39kOoW+IEg3RZl40lRiWZWHOH12bHlRE5zr
f0g7lpMsjv5kQYmG0pXJr424OGykf+DFa0t7B5B16stKd8Gh5ZvawpiIDFoVNAyerfIWWv0YGBHV
nCSbXN7j+dm+T//FLhsS8MXP3FxnDGtrXZDqdTjDHNgCv/73sJ+4zQyy1jlloJ0eHuScZa4dMRRF
+LCVIF83jd5dgthYqQGJiUzo7BHxU6oow8158qaaXQqAxg0+iMh4FJ5nag4TQRMcKz+yv8uZmm8Y
Vd3sPV7zDt0KUcClRwFxExbLKc7nj6xmpKl8Ff8NJ7GcHbTIyIQ+/jRp+eSS6F0TR4ytKg5QEd1X
BofFYNJ/SSa7oBALMeKPi9sN/pMZHEbOZRDt9fkVOcu6VxX6viYgOSKViaITznxpgqWiBphfVB8L
BeuH+aQzQFhBGauw7HzFWponb1fByDPIBmwv3LZuuA4Fh9PuLKktx1t+i0o0K0kZ/0rUEtWzDWzF
HrK37xnoeejiEJ+2rc/H2yFekpi6/NjCt7MRmaqhAOvdy4W0DvHXs1UA0xn2TT4PyA0sKDGgfI7A
zEunHpzf5RkSi60tLFANRxbKFrp92RGoXo472HfunvtS4a1IM9l2OX/H3RiBSI1czI2QGIR/UHo4
cQnsg7aww34so05Y48StxFki9mOgr+wQEihYCb3J50RTQJaUINTLnRXI83m5AgHQcd4WA9ugYMJG
k91aKg2UHf2+q32Lru4bqLhAPyElaUjzsZ9owEVXDUbzLBFakgNJ/CcMyo/ROkYrESmxQmDvxR1I
rIZ8w1SEqHNH5jT4l5JAjeFcmT1U6CV+my8W+G5LBQznQthhKstscmDFfBbqTOQi9CY3NNtKjsLA
056ybg56PyhCLaz7PbemQ1wHzVxhc8s8cepiBk5jkirhGDCzWL4Tpvy3+S6W3VlxG0lUDFi6dnD4
9GPFMNpYkGTm+zBDMBcqyYn45cTLrUhm5E5Oi5yro77oJdv6NImuO4kWsm7CGIEgRXrEsXfxdYoa
Ll756e5ttwJWcKUhaUJ7fEjlfQP7QqAoAJ1Ujxg8C8b2F2/CsSJrbj1kbHcotGfIcj3rYsvRrUQY
ACILpcix/luE+kc6UpIEU1h8ZQhQ6IyUdVXzGDA6Law5dsmB2M45abu0pInaYzutkMx6qXITh4h2
d/n9+GAAaoxCZnfdx52q9OV9kWTUQBftiFa2SYuLBcN9dG2Lk1XBy6Kww/w2k4YNuTcYV//E/O/e
Y5oYRET1fA7x/vHNOhcUbffvtfFTdg6luNxgbBis94BXgDbt1Ex38t6xxlGMYRqL0RuiU5Exuizc
k5ZXmTPSWn1MaHuZOF92UCdQSkh2RZrKU8xtLxErX+ucU5PX1U92ir7sZoAojEU0ssZcQ8YoK8d0
1oxCHxtegkn+OjAmfrQZ3P6n4/m6njwvwydZuWijCP7j0NhBb0fDGnpYFmqTwNGDwb2QsIpvYfZb
1HsDqBpvkMDM9HMf9beciEhwalmSs7JLaAkGA6h0yxXcV5Xq/4IU+w+fPnmZtm39WWvVTo0peyz+
wYeAQQIinTnJn2lo8tm15bzWz5ZWNghL1suUAIHUVP1L4kkrz7WwQRi2RM+8K3TGT+fmXVrxtBzV
/sl6DTB3ByVRCDZHp88utL2XezrV8gDA02jn9HpH+KOJp/HG45/k2C+CCBkzkzEMn0zX7qmLhJ5b
n36iVs6DM7pn08ucqUbxWevBYtStuMqJgQmXwfcixiccy+7kcL/H56RSo4M6FE2iZIem5HPpR42y
FkUQJrj/wbduWf8YSkvrOkXB9DNddLdFOntY/bJWjE3uvd9tbtG/anvKAnOUduclOdKkwS/B9+wx
KK/PEeFJohhx3O+DSBWgk71K/K4hM/dZbo7RqYuGF6G9Aq/rb7d7rlhs5ITeReKKA6C97VVk6Czt
WmzlnzI4hhhbSuaxkn2cU3+OIUaQCuA8yqTKVT1Zc1l6HCaCyvZrcIUYyT5V5mwf3e4rhtOne0KL
lspS/SVLBoSHUdVpQHjVdCbpVtu8OF4fndZcQHxEph8GBsX8fmN+E13dtL9JO5dcJUZQpdumeab7
j+EG1SQT1BNb6qteDsPuAR7IHfuegZ27j5XyEaaazKHd2dxHu907ZIlcwRmiUaGjKlx23biU3GD3
PcjCr0Mu7KZKGjCLNLPeiIMFjBJkD3Fu/OcwpzElncO5QYercJvs0DjOsmx3utr2ORQ4KxzdqNUG
9eQvd9OXCO7sDphnp8q+62ESsSYWXXtpE5N/xkgc8A/TveL9goUPPPfF9ilYZgJa+uyxoG5cKYFq
8ME/bwNzOCv8qAm9ZcM3m4+ZsXIp4/Pmp++Ss4gWIM/KtJli2cYeV6Z366o2vsbGenRPmQPpB1CI
5vCRVrfXO7wTOPL/PdMxU/UT0rPVpv+A49d1Xk1YWT0yC3bbgYVOb6y9GZD3sYthP+LH/WoxNgZg
aiCid8g5G8ZIm+O/zpgC10VKQLIgwIV80ldEfyMGzpdc3Slp9MD2JzV+XnDUTDq7ZCk961wVTdjK
o/yYsLPm9b9WsARFwPvRSoBKREuWmc+sK0HLDOWcviDvG87TuKdMgxhhymsUoWdlNXI3Kj9NuHLd
he6c7bFHSQkAByamzJvQV1NuwATWO94MO1Ihh9qATdaVH/VsXeXP5IzCHk+PUH/vwJQqWYHh6wq6
TG1LoIcXanA+DfU/KayLVZ+VBBiBexXrUnEwbPm45g6woYnj/vd2+yfhJeFTMez6dgLvVsZ0GSqJ
lj/rpbT+eG+vcTTmqq/FbRVBQ2gYejFyTBRRnTy3DOCAsY8MndvqU72IaamebEJjgFMcgNhZ7sth
Gl49W4NNdFJ3aUNtKzTZDyrfg4hBrTDwHA7yNOj3aQpSVF66fTeaS1gmzFuw8u6KN5gEfEDmu6oz
N0bOkayhlXskn69ok+icFsrq+X63HghXWDuc/M7BLuEcXMEDzkKWnXJ2iVakrTbr4xn1WClumVO7
E3qA8rmmNHRe9/8E/bU2mptsBoontNF22m9sDQgO+da5Jp9iXTWFBhuACy6HXVwcOVyUEPOGQb4r
RXPHQAL3emYTVUzriwllJlM7JUuYlxTh+Jf0AnBp9M6mKKHY+uhDXiFLiE2cEA3DBH5h25uEH3U7
CzSZGJyyZscWQRekjdECxMOTJ1T3/jb5pv07zuzMcvPV7PbIRzqfN2rESUkAROlR8fvcvPASVMzW
ryuYrFtdn6QaD2Wx2cbAJqC4GQpiuCrgy+Bs//59BTp87b6PV5fzC9igamF3HnC5/a8v2efmJR2q
yRAjPlbio2BIVi3Dn/pc0Clg7y/PsZy8yeVPcRilKZDfAzwnryUbfHXIs8IBbWi3sTCZOADGnZBd
KuBcpACpUu5XN5g6Hj0UXvXA0qbqbZH0ZBCPG4psTijnmbeWtx4ssgjxAXKC4Y/pYPhwqi4lox2g
A2Zwa0oOIUTMIich2RFZnv3Z+WJ1vpvTbjYG+m0TrDzayh5pW5RsdjQgsz3Wr+JQUN9pl2JrmifE
MZTenRM2AaT5bVgI6iBIZAOicd5xpQIfmJ0wI7rw8ljPP4DV7idDLrFNIbSbhVt9eaffxO+8X7RG
ECC6A02PiI9+2Tb2cYctOdKGjmJ8thQfu2s5ykEnPDLvXFbUZ9v6UmUnRJXoY8C/ielVBkhy48i9
mWIH+TrsLEsY1NPWdMm5/INi7nIcIb1jEo/IYxFBC25n5DKrp2AxsDmSs2jLKcSFWR7vNUjClySF
DgL1YRUPoJI4tUrk6eibpGW04IZJjS14JJZiSBb+9KC9H5tAXiCUqeTYvN7Ft73e941PzrUWZ3nb
ta+c0jz8fTrpeCarfJfgoGqchoniumxHPWgD2W02SypbqekqvqF0KAKvNDgaEn7MPySqGMh/BSVe
YbddCev30rTsVDVX3w+X6DDBhIdUy98MOvz5N/lDpPkelTH9be0EoiZocaQbfwSRDMXek1dTNnrn
Ck3ItaU+Te/fTizZqNtJC5UNvrJJUpyjvSEzc3UWdYHYLDN7CYPNzf231mQWH7pv8/cfePbObTDw
heQ76CkNBaCxPcKlBdCai0GaF9iaOj61LdQx8LxhMpQPm/dhPUJJH7L61lIbH/jAATJTzNysiZiB
ShLdoNWBQ/xRuY1MZP3Z0OoagAbYT2n3jHZS/JXElkl5SLhLWb0BdKSfpgqHsMRGTonvy/hubQ1b
dxl4si3jAKxHJJvGZ0loi0KMv/+C5FyeCglvSkFp8qLgqfvqYR1fh8QSr0IwL8XP3J0Meyt+R/j1
TuuqmHM7+iErEqGoOliknCQ5XHHFZvKShQKmGjqmkFG7Lzv2n27SzbDkzyYv3FJ6f2tSvLiMY9zo
CpqG1nwmXeroy8eTiwIcaxmraV5TV89V/tWWp9CNOy4e1MQTCiRDpfMqNrxD6Dmjj4bUR79VZcGO
9ZmgIUFwRtKtkQuCx63GCMUiT0GMk5xn658ZisqC/crJ6QUjR22t3VYrBJB+8Ci95ENlTgMogug2
30XIP0AexblG5jIRnG0T+V5W4owtKGTnxvMNy8necWiybnFqADZAKQL0rXFnLSCy9psRbVmOSSz6
EeaUH52dv8RNSYjmTixeqy2D3QX5WRl8YaZyye0RHOvSFKpGJekQ7/TdnNorZzCRRv4eNrkRz8x0
pUiukWZTteQ/pwgLW74J/81DM4Kb5GXZVu+Zytk29LZKyoACtIUGgWviHRkmjuSLNzFmT4Q5QvlT
f4IS8Gmw/Eaxm7KV9uuZ4WLLKHUhGs/QjxaLJ47Kyrk2vLOSqMTyHDasCcPAa86tkUL2coFRzU53
EjYE1KmXtg6dB/2CJd1vxL57Z+DEUCIyXW7nDI3id2dM3RULcEGTTrK79gIlx9DQgbr1KnIQJoM7
9HxGK+EPiYevbNvEq8gWf+4dCFEJeY1I0iCGFaE0PZZO/p91U+lQSFNsbj3XT2hfZM0qJxflyr2a
l5xyp+y7SJGaAipNgOsdnN77MkV7S39S1tbimE9d03pN7tJdLfvgsocEenCQQ89LPhRzCO8SZBIu
WKALbApcG5xIz783qVUVBh7hp1El7O1cJBGI0Dh8cPBcLSWFs6OgtrucHkmhOXyxZE6sftGAnfgg
560/eHTkyEAAKrEtQ+MKlKd/6jeePZcBparDpsyH7p3sqVpS3npp9ih+gM/fhjjqVesP7b1lrDG+
jFbrrDxkj2iaETKorq4Fetnefl/qtqhW6y/QA4Mf+uS/EPQfHqye7RNiNMdKVh3IMnx/VVeN07gA
/1AQzOzi7a1qbHxKFBklsCmOxl1sbvRM4YXTX2FVYh5/LKhBSzLwZTWpwH5pGbTrSIXrsYSR5TUv
SkrFMxznaPartHOKCMNG6Ts5F5Cz10MsFL/S5ZvuaPt2Sebm5bRINWzPZ9K0XIaXiiKZ914td19m
gng0J/skqqiBO3UTFdVQ857mLEL4l1Xt0Cc7y6DNW+3kTLzdrUVifWo/m7h2/K1jbYw2RvUTAzm8
6twJznqbuUSGvXj63sH8m2f9QTOl7eRJAEFfj1oZ82Yd6WsYkaNsHvZIglVVMPUaN+CsTlWfYboz
l1sa4Dk7Dt9acwxvumNSzxrcgeVMT11EKSfW+ZhfrSKV5STVWCuvAFklW8OQZ54Qm/JnYvGkJ8Ok
n1gSa7n70Gf+I7pEHxEg8EQIIqFbqLY+KYuVMETngBvagRF29xc8PVo0pLSWXM7JtspJCmdjwCjk
LuWJhOwbspV/Hs93dx7JyuZTJ7Hmveg8qyIFLIzEKqou54ThLqlw+tRduyL9f1eO1kIHYsABnql6
DuNsmC0+2eFTGGNWupikBMAFJM8fy3E3IwykSrXDyBRiFitzJxueiKjF4OeVb87PGedNTfup9TVO
IfM1WwI2mhKpKZDvAQjqkBT12ciytqHpT+v2qIyQ29HVK53zxncJvNLdDrFVzVsunCsLYCnhlxAH
ettmLRonDFhWYllqZnKk4qmE96QyLssYvDzyewIOgy/jxf9ZFO/pMet6hrU7v3U/t9A3XT1+tchT
mCup6iUUo5oVGK36QqpXZAy5D5uIggynmqIVCGK4Q+DwHZ1qEkr0YFTCAE23wYhOmRpRKskAzVcT
qmK6QMrDXf1puQvbwPyrFTjHEbD5innmWc6b+e3Ijnj83mzEbASnEo76kZuzlzLC7SKCN1zCNcin
RHypK5xXai68RAlrKwCBMd1XAq4VlL1/kCrGZVm+VdTHi9JXcE6tLLqu0Mzh/QZ5WlyL8paHeYTs
l6ESCDt5LwUPK2rZuKpOQ2vQn4PPGqFfcO/wc5vpH75nHAxtYVjj3t7wA779wYwCsDrP7PSnmDuS
z0ZZEaigDbFbra4Yk4N9DD2LG6s7rAkdqqMfNHFpXBBOeVRoayO05lIn407oKEFXiHVvFd/2DraY
Lksow52W1X8ylq0E+Fx1ISttQl1sfkJ2VCEoKtPGM427TcpHAgh5R00PF7An8YemXPgjkrnM87fq
NEctCNrRdZwpVylSuumgHskq4r8TEdN/M+Ku+kVSqdwqhLlOpbTciWYAnQncv4u+Gz3dlcALSd8r
d4bBS7tbIQiOsRYXEX+jXhqHG4vuETF0Oy0UkjiJrFCpgz5D0Mt1XSpTSOB+UPb9ngEjaiw1p2F+
7G/N1S3BzNLFjtrZnwnxHbXn3m7EBGPgTEeV4cZUreuNRScIer0LxDlCHfsZ9pAozV8A192atCo+
/JeEIywx+nuq+wlAXEvkOdlUt98bV6shooXPjbvvsonAdD86EKRwAVgtYTqTB74lB7Ebre6jChpH
5jVp3tFbhPmUyOcdpdLpiVjf48HvpYGE7XbxuvVnENVB89FcM1z4cZrOsWgHypwBw0PDoQkgdd3F
+zJcXmdHvc+8bcwK5SyMAxRskLF/IlGygDSgHtdAdWN6jpr11g9SFIrQhL4Vm6sholjwWk1mb0KO
9rhduGTiZRjXe2UAYU3CgHbJzaDo9PBe//EaxpLUZYBRiicIEIu9zVNWcJK3B7WurVYN2P87zLsG
x/76WAeYe3a7NREKxjlNr39aDX2KTsak5nzBuWDFw9ieHdavW65ccvU3IskkwI8xiUDkc31QD6bP
77sv1tHDwGbvYnV2Uy4EvfrtNHXLt5bNWP8gFAvohFeVkthrd4kmQe4X46nXoKcxxi+8S8uu3TP6
zYPht70gwwBBA3yf4PkDdlD0BKsiYyj0K/DZNPhfp2guaMHdEfmekZ9qdoxwOeIFHP9lm+dxFo5X
VcsfjdpUVnYbPBO/NgyZ7zoQMwHnskWk5g02CJhkMxWaVkmQBocUmGoHltfzTeD5/+9OOTehg03W
5A/+MVVc3t/od3+c9fGVL0sOvi5Zus5gmyHEg0nq1QUkMl6U47yuEeMesFjDrZ2xdl9NVMukir1I
YcbS5SB648lVmlz45LG7PIilPCafFmM9v0haShBGkCBRbjIUZD9vs0lfmZEUU7ZnhfydCJYJxJRO
0TPREjvpZBzb3Q5Vu5yrceMuG1ogwlq6L+kzG/AirF/dio3hPy7kENGBWKPx9SJnLdiX0cdjs3MA
+V32m8SZnehoewvxbnARGz32V7auTIqhgaUmvstIsjRy/jQXbX0As/NFk5N/eEpCoaYn3+iwA4zh
5y/JChqitXKFSH0L0LtspRZf9OKwrsqibGD2a1Nu6Jotx+IIWHRkHSVnEJ3tM7ck86mPyr70HPiZ
otfUcbPxtW+zfzwWuDLH1kk+ZI56gv/41/GJ+EM7o/DtRx5sgJ9Rh2nM02uRDIh1pToH4eFRmKio
Kxutm+Ua/nLDotHyBl9aB8l24YpKcbEwIy5N/Sfm5wHGZowPlDfHn/aW6HlZ0aFX4GyCL7n28mCf
yuqESEZZckMlOTd2rj1+7UuX8zQOzINzkherXxVORM/OfNSi1lmQl2wsYomRUVCE7dR7QxxKiPiD
fzruZuhxt27bozt1nUzScdXJLqScL8xQHCIfFg4O+gXfZVfnduiIYWCyZBchgVimQyG2/RQ2iq/x
1AEYyH17yfPGATFuj3p+vXc/brp6YhBifVNn2sdJjbeEha2LwvltbU9X3pFbS6JyrVPdbL3ssbd1
HpVU4K4thPHfzOnPELZXGJ/fM4eCsvobEQ1a0IaVH9MiBJmAOAxWj7niKJ+p9eL5n+Q35eNQkn7+
Gv4fTDqywUNOh2F8svgyiFjfLGjAhgU+/hZ1OpVnauX/KZ3KmtgH5ngUXjeTcRwjwnVRozzk3yH1
9sl4rTaYuHcvClox3Z41TyO9Ba+0eFF5uo7LLJ3wB/LzTIGslGtPHaojfZSQAzej+KQSe1FfFQwh
Un0RWJD0ecPMGPk9R7/T2Gj1bEgwWZhZDzNJefqQB5YtoSjzlDe55pwWozB4e5UV0J+LiaVXwYqe
immEpqwfTLhsd9k1CipwbmzP4NijAoarQa59rqfL+C8/ESQEjySgxcEhgcXAz5P0Q8zmbXEgzFMq
a2t4TWtsHfnPG1G/PikpwnxywIlYB1Up/qkzdRvVqWnTW1QlcDle5wHOm10x2tuqC4+UzPwBlZDJ
8LoLurrbKFSWrt9fUlAO5KFv/351SbjDWJkznkyTrkMPimHkAI1/glfRR2yyxmnGW6U9neBWKgmK
MFuMyXaH4IMcjqGMXrvfdcmau1qDI6f4rB8Moz4VAwKK42qbKZtfR6sVx5rly+Mfi0EDnax6BT4e
dCSJxU8LvuXviorlmz4Uku0xerMYPLbNKqSxA8rZq9XRO+dRKereZP8YnB7Jz8G1Nm7ZyzSxJm8Y
fi/zf3GmokWpySQBvw0Y+WJBwZ2XJn5jqh8X2YB2J1xNV6MaztqNNuQbJNlgH+eCWeGYwY9nc4dA
OLc0j2P5BFBbtEOjhm/xIDa2dsA5BCHKtUkC2FBp4yykTJTf6fyW4g3LtwLtt90/XaIsmT0LWgKP
NDnyrREKn8PpdwIWNJTI3+lBHVMWCZb3oYfNNKRcZT8yeJDWfsIMf9lW2NBI41N0XthU+X5izdZP
rgbGNCwVZZc+7pwSzVJS6+cXRFU0b9VpavvEls54hI3mt/utv6oPVDR4rGUYMv4yGDRKljTIJHok
klCgdxlJ+lfuYtv6eZBYRkHKksmeY66VAHU73Ls3foMEuVj0U4cFEVzocLwf21aYg56Ait2zZwhr
CRVrkqlYQccxplE+FbWd+SEjgzRSlqfzbdDfChOho//RXSA81xINpGTEwkdao9iwTY5S4apu1oby
v0zhJjtQ6nDlZJPT9BSSwK5uu62V4skzJfwtauZWGfhOoNV4CE5/RxbCcEOqGfkQJLCHSntytarq
GkV5EL5pyD2SYUxci1ou4Dt3RdK1c7wE3CA8iR0/WrfYqqZR+s/osEhW2Hz2J3ULiy4hUoKJtjh+
/KYEFrW42z6LXiLoka7P38HNZqFk/IbBC+0FsrdxHsgW4Bd6RDeHLaXKIRKhgiGZ5KE2xeIHrdCc
ig5fro4EYRx0M6i+RWTtpZB/9vUL37G7+jR+TtBXVjGQ/g54Ashjxv1ffV9z9Xq/qaGKqMZl5iqO
bGGz3j9ag+3CtnAw+3a1GOmPL6RHiyPmTwQHUccxTgMYQugkCvEUaz+/y251OAP4dpo00OjEyyED
iDryRlgWWUocCnaDNsxlANJTO4u5IAzAEL8sZK5PRB8MqWGS3S10u/wf6gsLmaRIg4FK8ekvYglx
8AGg/ARvqeNzhxdMwhzSPSzi27fFvfQWt+gb5njHHJ+N8gNV4muUuP/sme9V73NUWlj5MxlQdJ9u
Hiy9F+508BjhdiQnz/keztLtMVMQXUAm8TyUzwo5/DIXub3XZMZjq3UMonlceZH1GL4TvLD0NyF/
eG1QouEUBH31VqMVhdnIx1f1ptX1JkQusUeTSnygj+x8Nh7RhP1K0No6yvwfc405q2T+2WTzlvWO
27XRXggvoxXKl0mbJIJXnA/dHR4gUoyf1JBwxXSHcVI3rA0XDU3lhKWHb7hav0fbFE+znfaNj037
OAslatwwTs8XaBWTHKJSlPUner5xHg9BHBTYiMQiMNASPPH1/lKS2AUBPemKdzsx409FKPE0INvd
kZPmPD5w4vAhFEy5V9ruoea/uc/zsEAiFgVaRLa+8E5uHxuM4kypDfqELDa5ZLvx6cv01v0yB9xe
qQZz7VzSz/DtR7xQkcDLmDa3aQMJiB8ww7AYFFEnbqLFdSTBoy2XfFDMCsDYajor7Cy+v/vO+HUm
rxDpqbzIq12YRaOjiBKjpW0OFhGVJNflWMR+IDKNJCuD5UdSE+11VLZf+gFA0T4CnmNNXQlyaSN8
OyMRCdtcnFCrePdL9DqK6uJPaUvYvkey0YWF3jTAvB0I9X5y1oJLoQ4zXrcyFzPqo/5+h6qyCTK1
f/BqZMQAXfHJfaFQKse7UPuEN85I2QEuHuAI1I8QXbHzhZPfcvjXE6WBrDidKRbIg10njHIncIGB
J52kOwdbo6gHSE3+p6ErpLHr9EdNfzg5XYytL0kVp0wAJpN+wG299Iax1xRP7ZJtLwlb7dXEE9al
C75jJxtUVjRnETsstJsTOK8Mk3lzz8gorsuw1qg4Tn7RNZxVtNDzh/H/K0EmazLHM3jP2sjNW+3/
DrUnphHYqw0GrEdqkwJx4gglpSzrjVT8oRCpwPqbsV5pqlDXWDfKtQ1TyWBfZCbX4PvCzxoJMVVY
zI/Z1snkytkqvFaFlMMF4WgLi+DMn4Po0szYP3O7YPKYorhctg9x80Y5dp8cS0leYcR1BZbRBZf+
ZyuAuxY3bw1VPPmwgFiIyarTqL0KydWNMazra85xq14OuHllbWLFHmXtbKnLx+IUKKxolPjZ7Alx
HG9V/Y9aVAZLMyh719Xk0Ikl7NmMD1ONhYkZBMgSFYObmYptHjhhGXmBwF1DsIuXl99BChhu9FqG
GWs0Mbx7ONSUTbNQ9rNUou6YPdpwoHUROP2rq/LL7pdBfyBAPXa+BFeGVmtC4fcWOQbW0Vjx3JMv
RjAK+CFoNevPqFlpjhzlDKgOgmnb8iVOZp5DZuufbPfmlePt9Bc7BUkorWuOjY4GgEudjhUkHkyY
eM2dDmfDNnI+CL1cA7628HuVe8p5pLQmOicITCXamVZLvhQqTBX86f/hujJd3LdPvh535TfmCJl3
s1Pey196vVgQ7uGtxtOFYLONTYggwmSV8i29AaFBm+XsnadtMaGmMD4XDWCEdpFF2VBFQWS24yJA
K4JS7PmptDmK6ZuLansT5MMdUZMxi4FTT9dDdMhW7PRkBmSLTXEZHcmMroD+Q692P1oDKTLpAqVb
xh2S6CGOOiMpQMpczXxo9/e/T/8i8W6F2ROc7NqoWekOwRjYdYZjzLVDDEsBLa7jg+bJVqmJqZeH
u1+fy9zTWDisC+1WSNAgvPD/NTydlLrvoRZlcW9zN/Iqflendaqwk9aLQvvFKA7ReBdlONAQllTa
EczPS5sZSxCfp24vFnUKejykA2zFw+Tpl03i9rnrhcGw/KrolpHU3eG1WttZpYKR5LzfNmzAeTew
HXJxh+jcATOLTXKze8oRr43IjxyV+/yRv3KQuQwySrIz4ZsxotYYKg52bTsIDXzTZ1aw3AbnX4Pt
SRlqjr6CD5vHkSQD1w3UZthBdg4jqVpA+jrhGNHsr6m2IPpn3x6+gkOtPHFtCDjWS399rWs/Pre5
l9bl0Vh+O4DN80J9KZ5iSEYCtP7IN2FiivJfIFXymlzLRe9Eck9V4Z1Ds6HBaRCiAHrTUX3kp8tA
fvC0kYh3OB8DOZ+VNv+pTdq92HlTJ7QiH2h0xCHlKZxbUtMkXbQFxr/+j+PAvumTKBetA2fIZvYm
aO1xrIqYg+MC7Dci8MmwvEcdTJqu8VQX//+F6N3HI51zHPvu39q+Mxx9two5eElHFxP5Ol1H8Rzb
K/47/C5QPKHSk+YPziihiL7TPQISWuzbmQ5Dm07cNSziW08xwxn8fxeckJjjrBkiQlYi08flwkbF
PUzZP7nTFBA/L5kmVS1tLPW+ObSIdnqFETYlt0Pk9FmdOFE2c++AD6+1NLlh7zI6EehkEyDtomex
6F9eqz9Qz1zaXXe0tZIGFZzoUsfxxsV8/be/IahedMSVa85Au4nHESGR1wiV05AjoLOzFlrjJWkR
f0w6wN/mKusTvrKceqOSI3hxK//VoddzU2bmsVj0Tw+MgV8GoglqN4atjJm9sY8Nquc1BbvgKoUT
ekJ/bZ+yR9YbROuvM7F10k20DVNAXML5O0qmTxFesM2FTAhdHGm7CUVBaXlsQLM+V40lpnFDgtH2
NdYMwQCTAuo2NDkyFSj4+7D8RoU1tl8MlokhkiKaFSDFJVBJMWQlyc08LH3mal2T3NLCaJ3sYTtJ
Y7YejzvoZaNNhLerkpHTIKC7bEb219p45d4UVTZBvfBWoCBfQ8bIHQ1j4wIixhH1WY3c8gd7meFr
NlZhdw3ORuXxDkFtbWdWUZUQp9fC7MvFQFye0Zk+B/uo9m/M+oTLWU/weM4Qhwv3zJTot32xawvm
fQ0OIu+gOyZc7jB1VSoJDUmrq5h5gO9fXW7YttN3tsGS3QLcmfjEqwe/LXuSxH0E5LJGnLraQ+BG
LTPPXKIKPGmVlGyRS6b8WWCUjNIrT26unwM0t0t1+r+pLeDby74UaJ8eRPplcl8zcqC4fX5uQ+vA
0916UeYKcRUGXRu2UCy5Tz88hn1ypUEmbSI9f8RIQ8fFUkINH1vroz1n1StazXtKxof8lgtCQIY7
oAqmAxc/WlyQB5WcKNkFCFs1URBz++bJbKjT69ZpPrPkhYHPO9FifboEDVqMajX2qQNXwiiDT05l
dz4ixDcbeB0BeV/YkiKJ8tC7v/IFgqrngydVPQYdCcDyaAEhai2A4P4ilmv6RTgAG0hTszMFYXDb
dBzhcJGBjE3b5P7cmVpzaSAN+/lxVg4+meyCh5cz5ImxFOQV+PJpdB2Iw/X+jEXxNRRNd7YJcSZz
gZGT2+y4yrjvlFjfGm55jo7MEQkwY0n5KnYcxPRgNCQcAa/M21dVAbfT6mRO0coh2C2tM2ZmlkBb
w6g1uhtjsYeIfhn0h7TAw+Jd0yPr1cZVcWgBypN6SwUaNUnCU5sSy0bsFuigO9SVfHzMo6mgQfxg
LOdmeBp83t9WTLyzaR1LI/RhO60ULWfkmsjx91urEF1hwmxJXwvpPoZpM5ZEfCXFssrqeoyOXOvs
HZWwPCrGJjRT9NUBfxUrO7iKEIS28Qkxp9eBeeSQYlAbHYF2WgeY3KznoMEZg5fyG8u1KnkhlL0f
MQPaIp9YCxrwKtpJEs0U/2Dqp7FEIv98l1i8S+XO+xKYe0TDB/9jzG48xSTF1JzdoP6ekl8jz441
Sl+I2Jk8z2JJEFleZKkBqRIf0wzDPUTgrrCETGVL40ZwJdY33iyd3FksA5h8/KbpPsaNrwDnJngB
82vY3e+qYsoU8Hl0vLUZ+RqaQfktGhEFVenjJ0lpD1uR73T6RQKUS1VDPrubNXsHZ9MqUbYm2HvI
ak20FOmA+vlC3pKRRIPc8NQVct2MLfGwoZPYGHWqPMSJN5vug0pm9T3VhbYOHt4gfyz0KOk2m0D3
WCPyr1XUoxfoY4CPOA9+u8IShxej0+3vZNKzlg7kBqBYaqpiDwiyD6VCoCezLb3uSs2SayfJc8Fh
Fwa1WoaZnmX4vyMCfIYmAS28RwNd0V/yYXV8h5ZuyUO5cKVcLL9nMwAgMloehCeDtfGkKCEGgi7R
OvX8auZhfsSor+lTv07QTF7NKgjtc3A5dnR+kEqgEIg/BnHehY04sHIToVNZUVChoOMYbboDqJXh
xAOw0hyDmB6Kcf6tizo2s0n1ZSOKXS/sfbSUOGZp13ipNfc+hEf5ylJtnKT/PL5CeBIvJ2sjx8QQ
3r9jaRLZPjEfVg/Xp3wHWw/K4yTiQY6SWfmfDHCNFOcHrTA0LDEm6hqKPLwjILcuPvrp7Hfi0O7k
NClmMe0FlAlSCS+6zedgKHLv5Ltx15+/bS4XXZH2YShVoMVJcJKzGa11HdwTUxWJiCeyxqPQTXBE
jw09VjiXIVvrbeBJdLEOT+K/z4Gh4TEY3WaxObjPKIOoLLAGW8/Tk/1BewB6Z6QyTTWy2F1hkEZa
cnd2AwGHdTzAlysJLdqE0QvThnjmpvRx0zK29WdJcuJhPVX9AdWSVdKvepWKY+IRDzBV7pPCK//L
aN6C7BOvaXxtBluXy6xC70oNMLWgYN/tpu244vp0XGCRKyn0h+TeNuZwckHGEeQ/Nwqrmr6mjfqf
accgOs3aUGD6lsjdtEn1jPGn+EA7SP5NAuW9FzChEuWn+fzRWddqxL51XPBLFJuI0zoqGywG9o49
8ravXXnNhQPawTKH+KTbeDzDjwxjFB+fsPt4pJBRspOD4z9Azi/Vqq5r4HQ3w8O/Ha9UOhXmr8OT
spC+qo4+ueqMrZrcNbd/kjjOIK6pL688PCvzvOUdSOQAEZerhlGWH3e5kAuoSr1J526h5EoM9i9M
nwRc7VqeQVocACr9v40S/Ij4K8FleKJlfm+UfpkQhpDUUs+G1xq4UbP8rfRQ0Yghi7tu0kaeCD3e
csjYHKRHoC1Usy+sS6wHDgucSiCmeOqHhY9/L+RtftwYQ/ZLJhpJ9q3Vq203RmU8vhD6VD3bwiGa
EtHw3j00sZrcKX0RBep8o7lc1iSYkY9Ahta6hpfg1x7ma4z/mo9YVXQTjgd7nCQ7NXuKsTIdihao
2KFgaPDbPpzKKt0hphGFzrahhH2BVKyu4J6U+GAqYwoZXXrUgDisZompYlFWu4TQqkTaWEpIrSXg
5DDk5E2dN6uzPw/F46hPhGH6HsagTB1/rddpO40p+jOTSB8okae3MrKggPUjEu97Ix1Mk8mk2fvg
IRwJlrFMT9lBVzZ5q+FlcCl4W19Z4JAocnwM0nr2MOzmCOhxCgwjPqIWa3fSomIy4FNhlyDkPwpA
PgZ24wzbUvOj6XvFJB6h9DBXyb48C4ZFDYkBoA+so4J6AuImmTWer2swFM3BuVe6yaAlMES4N/UL
bJpC5T8xxjfeEK1LtbI48PZ3gRkz3ktQQ3f5a1YGoQ2OeXIG62XqAkshHA9frMm7ujw2CLoT9yqq
tG/xlWRpzXw4brff2D7i7v4BKo7j1RsuG9KoJp8oRsoZTqjJxn2jDsdJ7DOQht6ZXGeF09wMIfDn
tRIOhFtIUZV675quUxv7xNFlARV6nMVGMUqBtYZ2J087sgKJ1NSbjroI+HvR0PO980t2R660zDDE
fxU5ks2kshq+Ol4oLuBWSpi7/1K03ZKBvaaG4m1Hd2kYLvRzbb94s7PAekCM7AkuauFZL/7SWay1
5ZZk7tTOqf7IjVAwkA5kWVf5EuPpEyv4H9tzQ09bloeIlNSP6fPFPEvcyQEtyo/WbM1oX1Ilo1T0
Jg8Hjc19ZZia49vr+lI7wDt+eWyfUPqPlaOQbn3fVRwgrQTgdcVFUTXEb7SeYh21kZpo3ixqJfY9
0cC6afUoj0I8yHIOhRxEMuSMSUsToZLldI84PDZoleVwWYSL3ZKFohFuMsSvGhQ76G1MnnSAF+8O
28HXc952ixXRKVT7aVOL+tsGyAuy65Mql+oXOGSvySnNcZ7WQg5ipD139hVHT952s9DuhNcTTWjA
Ej035G7RrrvBrotEqTvSVGt/9O7De49aLjveFGeGKCdVDLQX6qV+T2D5oWX8tHuZI+r1CGucjXHw
x3nLm3qYYXYYDxUgWvYRYg0pD0fOpiilWOakXGae5IdAMie22cd3MIoiQtIZ4D438i5t+m+XTD1D
elOCqkEOmkqs7LzGVwmZNOqxS+zYk6CV4rFjla2ULt68x3Pg5g9KVGoUvMkLq5KZBHaSL8rFuXvO
/XDP6BgBjhkQ4Grr3FCeNmv2SYGRr5B205shl00YmdA5Y+lLXD1uQFY93ll25F8H7xQ3ReqK63Xw
5SpkdXAjR6nBsndjLUSq0A3qxjJNTtvLI2RTOc1tSKvY4FYwFf0555rFekaLy1OKGIdvecja1ihP
7HFLsNFk2ZL98t8D5XYdhkl6aG3RscPnDw8dSosXYzxlBBk40/DuLh1aL99KY5J8LbOVP0cOg25M
YxDLNScqVbSPx41qHOOneqeKDeDFHUXlgT9WjAW/j50UJf/sHv0CHHyD7k5cuFC09UpzIqMZl7e4
aQffVTCMmChzg+csNFAnQ9SkfTvEjVQU8dQycdkKp7wKjPvdGeH2ECYEl3PTKSmXk+32YMKnrcs/
bs8W0gJZPpeAnr3jZyesF1gsnCIbMkdPXUk0xaaYAOf+thLzxX8RBm0LycESJpn6QK2zGnSNmsad
NcKzrDwuRXo+rnUn1pG75qBg/tKrV9WkgXQXgHXeR71z6/uzWEgz8KrFOd/mSZN8CyCAPhUlw+Wv
zKF2oRVx7l8VBlMze4it2nR/YC86z79azrbi8A02rS5LOTAbWSlN4Rmd/6oROxuoDJbfi+m5+LIS
pAyhcM6ZUZUnfbr0PBqedsubOR6qUlx7V4XoXjqrsrvYkRN9MF9Jxplv27UHPghMFprno3P5tdGN
zXORjnQel6TW7p3u73oWcNZJhW3cd4NjPQXwtvAqcC7SMpL5Gvr00ULLX8+9iO42SoFGGfdEUpzZ
aLEg33DhRPIRlo8Z053A/GK8DAcq0gm0M+NjF8TlHwqdt2dPIeOVmQUFS3C4L3rn4Xhxxx3Ko8ay
Iv6/hYQl31PZp4rlOPqrZnCwtT/GqPUDxx/BWfHTWvmsuXBXFXYuAyyDoaZcVbKr7syvCOD79CL4
geGz8KUGtdSjIAH0SrXxAN5QgG49F35c5tHPD6bdihZ/6qDLmlH9cdf2OOAmuDVw5YP6vL8fq7zM
QLhX13hfl48gD68M+eTHvbeB6jWZ/AJq+4+dik1gyfyHDC50ZMRAQi7jsgckUM6zw98DR505MfmI
Z7HebFafUhTE4cvpE/oQRJPFeqTMhCfow75Ir6dW1QW1zlHMLZhq66YQvVkWFsPWiRQGyFpkpMak
6Lnd/EmSjBIFGSEpaMHkliM9Cw8AJ754+Av0eai6TKUwgY+D/PKKGr45MVdWEzn3Q7spVw+XoqJY
QgxALECNxvLCKsE7OMzz2WTkUMO5aG4DIwTPAVqzcq3Gw0zTuooJB2xBACLNAKWivL3XcinKBeul
sjIj7uZo4Yp6+tIZmoyoC8G+JIj+OWZW7mYv6lhSVry4IEfkxJ5471g3IVoEyf+5BmwCarjNSVio
VPi+bJ9My6OkhKgATiMZzvhSbP9ot7L95hpG3F2gsiXbsuhXMKu2pLFujxRMeX/tr5II1T/VEBY2
lon0PZ8+x0ihj49AxJLUclwK81NPptUkdCJwEMZs0DtMD9NVHaROWBUyYgzL1gtDjt8kdHUk/c2+
o3j6EJGJUHSqtxOcwlcj2zFhO72mBTyWIfCLEzYPW+CBo421ePUQcfQkzJ9V6octJslRfRe83h5I
n5mb7BR3CC7TUEKsqTT1iRgsCaUbOOPtuHm+Ub2dH7MRh92mAj4g4K+UIUmymJNe1lWclDj9gMIA
4hCmFECAGgcx8GTXrPtf0n8nKsmO+nNn+njQZRDK7XmxclIl7Ip26eVCTHYOiZt+4uVWM+IMbP4x
gohF7uQ1kzemBw08+EeV3hvZHm3UgHDU575KjCbCtmonY+qM0c7D9XL4x9ZAn4izGgkpfIVrvhb3
WIMBixfN5dgeDI8ijAweULoniN5kL8sROTahp2PvSEOHkg9sFzWyihSMlJfMg69a9pT1yD+GINQf
hbYN4qbx5uqjMk8S9FfAZuu39OtAIiewi0yYO9Zuu3qwQk5Y0e9tpR3f80pqeWpL3aqP6neuzLY9
O1qTqwOxHy2Q3PmpEBQL2TmKXSVGuM4JpSbHIrY7f9s7D2e+C+xQ/SsOCsZQNldSqMuaIFBka0hD
QxwXk8U7+Ar8YX/ewCXK2Dp4DjlbQF860pLwBcMdDbdXmyHSwCDBU0lKPtXHB0fg1tAdkyk6nfJ3
mIpPz98L8+Y7C5JvlQevUQbaWMVSOOQlxqys7JPPQTrLiAk4VN2KHH32awwIYPVwBdvhPRZld6oZ
/2DCRC8/JRNXX/Azdqy/aRKdX1bP/vrdO8lRfg0i0ag0vnTkxfX683gz2IIzmt3w5witzkcTMT+v
OsCLggBTlsvyu1Pfa7F/Ns9tnuOrG79IOaMoQXhkl19eI1gAgzxs3ixhrhnxl5CfYWrjeY3zoVa0
8SkzT+O/s0+yUZQlnquCuVZrkYmWdjfZNHrKXrkh73Ouz9x93uUmIXCisp9sN2k6Ny8CISfM35Nj
mU9/5SFZMJaSfWQCJO86+tYgX/3TJbwaOIT8BognilP2+k6071X99W5tVarDdZqx0EBNXYpC3+OH
T3/oiaIVbNhAJkEqDvCt/ieKMLGiemaUbPuaDsEM+plhPRVjD0vQ2ngBrOobicTQJKuoh8cXGolf
ZusVlKwE/nzRgPSbwguY4/tNSndWdooMY7B917x3rYf3n/u8WctjrIHDOIy2cRjlU70biZxPDD1+
dn1nyJQvD/6ZTBvsTnIbRIc3TOXmTbBTvZD6FtaMfh7Ixtt/g/W0b/r5vQtH17O9s4QRfTjX+lWv
vinDU7u+4X4WBmbh+An88+baFoSqPy0dFm9DSdvgqwst02k6mdiGlJXV5dTmC0XmE4SPmFqkde9o
b7+s3h1dky6RyjDI4WrnPqisAn74jx2vwsyY95S7RI7lMyUNonwHhB6/R4mqOsYB0HvdkgL78Kab
iM4AR7pz0tHYjXMh0y08lA7l96ltWU2GGMhL8O8uh9HLsyvSRq9/3RpoTzIjzCryNiKG9uPaFDtd
wLMm1RRHto8CkBGjakiAvfMK0HtBQRKoBaxKNBTBTqAjLDMIFeWgKj6uINXocjfTCZtovS0TeQLJ
CaXsAgTK/2CqYuOf5bQ24MWDS87TSzQZ6fnMkOiy8xgwxWvr+R8/gTBIUqvWuvecGFdnTSnf2rss
4KJwT4eAzYYdYXsdWc/UG8jciUgqfM10oK/kBv7PmBnizDQBcQ4mRP5iJPkO9CYYuilzKgNdF1Tv
oVonhx1XODQ6xxAMxYv0G9GJk7yo+vRhdDzVVf6CnRbqSmC7H5CcuFeocZ82dKO8INePYfsrY/nQ
Vjvyz/lgQr9tb00lfH3OeDrPyzKQS3Npc2v9A9ITvwuY4TM/V1UoCM0btb+A+acZfF0XmvMiUyDi
x5PX7cNq0V7rMlV8XXSCXIoLWu3FuUBLIld8pQKo7GEnuJvGi2YX96o8nzBSa9C2WcCLqaVNdcU6
C6mPXHx2ATwQWtIfvjqtZrahtyVOjIKLxAKU0n5ofxxCbBo9rQAVj0NVtwJODwT4wvDf0V0HmABl
z8U7ArfRZy3ndhAeIo2IfkKfh9+RwWqhoKquHP/4yL8Xaac/M/J4ysIH1E+cwFYbSgxBRcQJwWsj
bSU48/GMA4S0I8ze7jk+w64TDUj5+rHblEiwguEqKasGxkeKUj56DuMRJzUDTzhd4emGTyi69LFa
8vgG0Kp5KMmGioL57aGEwPO92UjtZZfTh3hveAeGuupRDvy5KJc+mpBo8IElww4CQQu45qYyzXT6
6BEZj8nvSpTKlqVSMeBX0oB0kj6Tfx0W9eOlmjQp70nCOEEvHrXPIDlgW/cIdLKtPXylbCR8PEzM
/nUF0yA4nu6yRvFEBtPSavb2gl8+Mor80P+dTXQu6tb8JMkHehiJkzDidARVojY7avGGTPc+3NTW
5V3am63e3JUY/1awxAXN1r+50G4iLtlLmqh8VFeq3COgMN/M9ImfDp8uNPnxqepZo0kZKZGt9gtf
jbBi6cRthNZs3VBpQzYMp2rMTv/Wt2nPAk1EWLMkjI/4wOMd85RZDOl4gqJoa8gxM03ZU+84+kGI
sVLU8Ic1SMYbJ931Auwm2TRa2lPvw3nlXLi21Tnmqk0XbCJktbkAg9w22oa2sie0f+cl8DTqQx1j
8e+6CQGO+z0J/ibEM2KarGD8vs3fVmAbhEg5GkC6ZCfxX/rsGy8ZyaFhlPC+cEd/zTTzFpZBcdQP
9iwbNGaKeCcbro3vd0c778LmC0aEjyBM0laRStehMr+o5L++Jf5PzQMaubskp4PPBipiTJpMGYuI
ENI8ZCZdf7YH9meCgYvpnLjqoeL02m8SSkJPgARhcqF1uHywA8RXzRpN2H9V15jJbuCxHKqyS79Z
pR3+r7QxKrJQEpAczw7B1lWeGxXQiemZeG82Ab6PxFX9UiCxgsXzU1+44m7qAzVPwwKX58rlEtnf
si4E2YrO1teWOpFcXdNxl3AqZ5NLxFzcPo7LYLgCSL5nm3RWTdQmwsEjDFvBflks06mbl7YR7rK4
+RuojTnncOt/bnLC2lgSjVcmx/CAoi2X5gwEn6YMd4tMlKAh47bV8gVobJ2xUT5UBvjowzXS0fRN
GlG8WpGCCpTORfATuEm644lQ7s3ffUxmNjVAwmJ0kPHezoEyLYdfejuuDNYIuAJujAm9Xj36Q/pz
CtxU09+6ikewpZDxsWCZTW+xnUbycuDKH65SDoWNwrb7iRjHTh/YfxmRNnmhUagSPOrAmnFqVukx
zg+d70+22QMCULbEJjGieQqhRme+3gV1jZCV2fEnP4DBS00RxT+5Fq3SlzBYK7dDI4vCrr55aCBO
0D/JHWw4GT2Hg+BcvdK6KC9vIhbUOR2F1+stFp/FFXtmVUrMpbJkYkofXo5yzkZB/7eiWB84Sh3E
b6ney7h4hfH4mZkQZDowzVN9Ck+7kW6sC3M5xe74UWZAdIwB+bE6Yggl/b5y7c/0Fqhnwx/PEgGM
BrqrslFTRpucjMW10Z5Su6NFN/t5iLGRUvG0VnubwXKMRwYff8NEJTen0t1Hkvrrv9rJ3s/Qpgmm
3cI+/4tXgi0e91RlEIQH4QV27PtmnuAF0TdBDi2lbmIB7PzgyXUPw/SDhtv9ocs46ngXZMQhvlM3
JDWoMbk7nL6bv5opRnYVQsPSbM3KTHiBJjizSodvMP7UM/u9oK1lg++gfWruoycWzypNrdDWaPOK
Cq2kBnRIpUY66a+yvhxunWVn0kWKDlpTJWCSCMO9FdAil+D+dxJFh5kePqRBLPir9KB0G5tOF7l3
vyLgQQBxz5IW9X3x/EcyACX+1XG+mJ6Y3LedFUk2aTB2savWjkl6M2jRHwJbl2LAOdX4f59051HQ
GoCq37yo8bFDVwoFZvUJyARVqi+w0wJB27zwdrRn7VYho9greR8uj+V3w3X/Em15IwiUqkDwoRB+
zZkSbCgOAO7BMdhjSnrupeCFYK3ReBK3jiVP02zdcTh8I0/S24/0bBnzEWH3oVI1FOyTXXIeku84
v0CrVOPP+qaWNTkh1o1No+8VX5N2Qsfvqivy2/iKhrbvDsU9FHf7zpsHOtI0VB5Aw4xCyJqGboO2
128vsVs11sE+c/2rYB7s1gADOpeo4iICFdQ6H70ffhXFKDrV4CaNvvnRToYSqc7/7QF7G/YJkjLs
J6HURH9YLU2hjzT+SgqukbYVnVv+Mb/MehltUuHNKY4gM/6ZcFTmckgUoHIPo1TSoOLCI0UKeNF+
Zvm7kIBqKII7ZE57Vq602x20DFwCaVlPV+kEN0F3dSeIijnCfYUGBYa2YApqU4otkDoFrhnEp6QF
gaSHU+0KGZ9cRd5ndO7CBFesiwHMTEpvHwq7Vq1hRuJm05bzTO2WKiTb/sfeaTvqlAo+Ntv9CFtw
mSEKd5WRwxqME7FwsvRaePo/UmdSAVmqnrUpEVEiHXp62hQRNEuDRIaIyQu0OiLMEOeGDE8iajyQ
mQWng42N8T/UPBeP9XG4wWn99wi+GeSXOPsBop3P+kIrusRWF50V0E6qiMxtjUqojEmPKiffNfoZ
wLSA3QgKlzvmfjgqE7Zt0faasZw/ZbvOsrZrlnk4YLmFO+dI3Ff0xAVRAYUkAq3aMOAmBLZgcFaR
ZbBN1kck0JhHnt9AJQ96QFIJfNJjetn0MBNAZCx9wQZMQtxeWxVdx6/R/EPMhc2Qahk7VyA0LHoP
lMYlCoOrgLlnux2tunPu4rNXSbzaCM4dxcGYCaBNPkzt/pvkbCgtmQjZ9Ld3FjHOzUTsLCb/8Vhy
kijpypnDjla1rDTGy8y7O0kw0gGH/NGgZfJu3rqrQpRI6vpbzrnzhth5MHq49U3LzNemD0tTr4nW
5zcdSGGt37vCNxK9pfWXU3pGEpoM45YcVGVtThCqQArVu3HmxX1FK9k124JZvyVuXz9fH2O995gG
NhvkImzskG+RqloFiDyvxKj11JoWxrXq5fqef5mWon8IU6xSM+vlhEALVPyUZ76ZF8r7YSZVIAX2
PXFWBhMZ7tOLtHN4b3VN8qt+QssoPZc68O9Ps2qDKGK7u1C7YRtXpf8Lsfj4oULAE+bllR/vEqux
FTS90ECTdENkrEFEKYCC7OjYaIO/4gr2oVp1dKrExbadugldh2E570cyaWnXy5xcZq0BdEn65POw
ymu7S8duk2o4ZqpK/pr5WwxqK+siCgVSFGGNPqjUEOwZhbWzzwMQrlfKCx1A/9xpPtvIxzyPAO18
fPCOOdRef+UG2mGaYga/wnVMQEH/zf7YTbEpFx2xIaAC+QtvirGNOcbA9BzZxZRaO12xtQqXng4k
CRsHdGYmVPr6XcHJNWYDkXwPsJMb41kahsbiD1jSzWaOlMlNB2SVfOluT3fU034XiFgioIGXuOth
wnkVY8UuA4toPm3qxugmSpoHgURzlvQ/dHHFVqvggiq9uoPp5hsjkEjQwQjq5jzlQ5kpekyEh3Cz
rFm99Hl3WVfXL+f998X4FhWVPu72IzCUpBM0XCiaG+UMuPcuTBbL+dg7rGDkPDUMDzFbGuGNCv9g
B2qplf0PxhlSbbKagdtYHTl0GdDHr80XKSCLeYCCSfFYpW7GIbxAH7V7QZlrrZAbDOe1l0soHw8P
3VjgFEmOz9lYr35oi4u/3QcnvqvcbIaEjXJ0gXm3bokvryroHtzjIZG49F0zuGZszZmsfH2clczu
m4Lg9X8m8j5EoGwYlmlgfiicA9jh5s5ZoB/UPEMKqfZmcfY7+iPwNUf5QIEuPWYXe+JKJX2FmjMj
9Z9MNbr+qG7hT3VUCAzP+yrgLjKn2Z+5a9MVMJjVdgrK3edIgwo51CghxToSmRQ7uba+6RSmDQ1F
baHI1hINsthl+PQdyinEdRNFrUI6LsC1HNAdNE9ZQglYWyhKGNvCpWjfNMwtiR1uBKQZOLPlW+lp
KTIMaya235U0U+qW/43qALa7U2jov/oy+kd6oN7wTtFCaVwArl/rSYrzakTcSdICe6JQlesHvRyM
eTusmAq4f78De/gigsWpoEb1KAnZHTU5wrBqA0aL/ROecEn8uOTB+zXNQC2f0HFTt5TDY7lZCPNW
EMtjJskPkmvixzbcyJR8XCZfFtqBb/S8eodBpC2rKfMWwlWY9cFKZkYBD0NBsRVhscgN3D5mZRPq
zQHkgd58CfZsSbfFipccc4SnABLlrF2ixFiIyZBVqd3hONEq8mAB6KUJu4asepb6NDVh9HrdfgFv
lt4NwrfB7XWexhikEHt2fGC+lr+RetCfLAPryuuwbI0KqWyAT3JLG+uo3q/MrcOwwHWEvDtFpzmC
/zxAhB7fs8PPqRK+llYBh8PNHUPT1x9EZJ0hLx/VG1dpWGwcDA35gJtnA7SfQe1Sy8Pewk+HTX8G
reAvlc2uo1aPUyo5SE60kHiMgWUYOTSjKG9yBof+Ji8nVIKhAIlpgGpkA7ScUSYSnNvYW6EUsc1s
6sDfD7rbCfi6nrs/RTR17soWE8iVau2YpSVKdUb+23ud5OTm56kLS9/Zm1/nLqxgvFdJPgIgRVH4
XYuPYN3JKgpyTcg2d74ehHSWXitzpgr5F4DfTAmdAyHuEr6J1zGpSbEHaw/Z+62UJimeigx/yVsn
8W+DuGFyhQlPe6EA/7yWkshw1lxIkuvu8rXZjy0nBXJA5JHg8R5xF1HWdw2DW74UEH1UtoLfCj1k
KbyDqmOosN28ImmE1WoF5YkQA/1Q8SajlP7EhItzGBpM6bfyZn3fnQXBPJzmSAEWZ8P1r6F+XnAN
k/DJNbpypubaVGbng130TxA6i9/5F7OKBygpMyJ6ZgyMvcFuNcxvFN1YTJWD/AoCM09x3t0l3QwV
Q2igk9tR9eB+Vqe5bIaRN8xOQvQYyyd8rIwP6MdE+vjCIqmnp/X0znfIwwdqHZKhbI1b4XA/c5z1
OqvypQ2gu3KhoDIMLwYaL9AxqQXMecvxkJeGWkKF7rTqLoTU4dVLvdabo5DKQUafRq8rh95I1MaA
mXyhsAYfzl773kHkAvZVoQNPXOdlrTZhOj7oPhEKV2TNVM8501LrPny668frvl7AvAKdcD3EFbD+
+etdcVaZRR0MzLCJTW09DNKF81dPgK1AbgnBaHuSbmWaMo93CWZPvZO+bklGdopu5WU0HdUdAF7m
dm12UwDtEjCnj/4Hhj4Grlhp4RNZA/MnNdWAKL6wsM3XYbyR0G3ynB6v1LL4q7f76TsRH+uKLCIh
vp8hubKtSOm8pb5mmMR6JX48JAbhwQzxtUBYeh9VJAEOMnhBkRlknBWeWZa0RyffPR62D/OjAo2V
eDqjlRdRKkXtdlBY9tA08QC+t5NDJdkINi2oHIbPcPiC7GXDdbg7DqKkBWY7fXEwXLMZKtnE8i7+
k1gnQ/GWyKILVtzi+qhpuEgTETQSWb8i7WG5rsEXLGZgi2De4GqPHhzi6hxDRo+8Z4eY01Gy7c0u
+i1Z1V9Nd02O8b7U9MdiQJ1FsNeiCuANvWNMXToks4IPeW/Nc6dr0F5O7/YvimYd0GS8gk2jdi8I
KGDQ6Bo3yBxPq0w26YMF434ZycdPLn0x4f65KstiQI4IxuEvmHmSC/g/ofVk5dKeKFuIocggTIqA
ZVtXp9QZtBOsce3OdOdR3YxMdurY4THJftWoxVV7PEwFjkWBzULD/PrA+CDOCTxgdSerkS2Iq6z2
DSFS7jcpvfAHDqXKtIM3FXiXa9n1HSnwMPsC5zJg1Hk32vY8eVD4KrwWl9YBKEcf7tOAV1FfID+v
8OQIMJBCx0jZpcMkvWQM5bFoE4DSQWnYP9ZqSJHcYT0mpVFD0+KLHwvwVVjGbKqw4+9E6GljqIir
DwnErRLiQ+2lhDbmPf8r7dh52ZpLTTrJKOY8LVaOIbwh4UwAoiIHPc2Qa/WttdwAKPiXlVb6ppny
Hya18zHxVGEUM8EBiAscnonrVwD8v4QpAWAifNWmmz9pltH3E6IYFhxYSsML6Oqy5wbFZabR/Kyu
dir5bGUUw/U6sqTwHvQE03hAzIbr8AUnj1uEFKv/ko1P4EtqLrbJOb/T+CDRq5WXnelvW53DGPaO
f8JHET2teXXwgZSl4FI1XIpAU48obWqOsJfjYlHshJtg0fVfAENoVPm+BfrdP4x/11T3CMjcyiJN
ybu5NEVedU5hqpEomUKUPvz2/Ttd3HiQ8UkWjrJL7SOc87NjfMRiETs0Cj6qevpklUS0n893vUai
fzj5XLoyf7ScLgClHZWjAvQvdF3/9dmfbmmoF71RK2qqX5LMQUO6OWQgy0EX8/+RT3AKdqfVNVKn
VCskCIB2LWpRBoOFUoi8qQ5ArxHizJkkNoktBdh8Ep75B20CBpJasTcQY/3LyrXTtGwC62VQIGv0
UgNY6AVz33tNOnVfFAeCOse/aKIToP5cAukZxoJK+aa+GAgQU8qhQ8sa95tlLo0bNngLDOPKDYlN
IPlHYIZ4TWSluqHC9VfR9cqnOxbLYxBL8TQPy/3v9P4DYXrjFZCAiXlgyKUpPSE/IUz66JPaqUCw
uH3qKbPfsW4dAZtogpozXdXYKn5JHJXhZveUbbieoAdrRoMwH35UWkm0zdbZyJnDzNTvhqrEsOnc
bRSU3A+K8OMgb+WKxOxGFq8taPnD0N4PLYqPJSXzMMF++1Ju8jFL9SBizUmhSMPID8DW5W2NaGt8
ZOe2KixVbIcjNX4IMfb1pQ0hYG1Wmf5QxquxfBHZWPcP73VtwwnKXdWbZ7BTfuW+fTADFhmSqh6S
7FZ9Ncb9Cxb6NSZlGotAPrvZxw5TdLZzzr00RW3RfMXTrFLVWeXK4xgPbQrE79gE2ZePxsTSKd5s
WXEUoKp9heUszJpjM2VomfYI2r9ooge6hwRV4dvYb9xku3E6uawv0jlfxG7ef5V9G5apI3JO52fR
JY2vl2HGP7M0RFGkVirh3RsZ56Lz/TLCDlmcv1HKwdvKcO7TnrrDhfsozvcP/AcWRuCGcK/MvQ77
zULyDWewRfZpBnRfseLWgH+n183ZIoYbzr02RXEiaK9RTEnqXJWkuW6nJwVCKtHjIbxFeS8GBRWC
z2yS4ehMGzJbOk9GJ9/IcRLC2Pnv6YzPeMfgLp+ufraMt+su2TKkNJJBVaArnZZmQjll0A/lRNt7
7uYFtBBLg5ALtLkORrrX6n0utzKV/pViyrR1H7IRxNIu42opleGe+VmKzTGTtT110zFwhbE/GsVM
/p2s5UTobpjTI4jo+Gl1ZcTj2fiziINZqMbRcZo1kZTt1RQC8eUvbCVJhYNapX0hkfV0IDpNrPLN
QN2iUNN5FFIIZ9eA5ciJ6UsWDGII4DWdj9JycAqle1LoOwJJwMtm/lCHINAejYQQ1NXSqZ76dklN
9z65A2aN8Fp1WKiXVhmF//rKkIUQvkL6M7H6KpAhEXnwYr94gfqv4NfaLEs0fxbgc0p9bo8CnPx/
Pg+ivItvW1ZMzHmstkoMXoTFuWZc9LBOIQmETAVZ6DrsVeSK4E7HK8I6G7viufn4F7wsUQ7wnGVQ
exF7MY8gcPasac+4yo05pE7TGZBsF2GzbHdTvR+fwaEaFjvwU75eXIkeEuF/sC1O1y9ahhEDwB3X
YIK+o+ltjA50aE9gvPAaQneQQzOj93hl+DXFolaKzdsOPyGSSwW/6QaK7pa9eZspjnGYabusz7bt
jBZ51Bf236CoAmSNh2pOqv1jmIXMcdPmD1GBmKP9jXNHitTc+1gYGNV6IJVLhHYw9Box7y2CNQpf
R3bQT01lFnhjVHvTk79iLUa6gU9ocTlUHMH92mOS8oE6/9xoUZGojY2OlQWS0tEQnLXTM9VnTM2A
fMjDTLT4YVvJtBOqSHS5rrWH/3yP4qI2KoVmKdMdvgC1Va2eeDIa30/NvQrcmhhuXK1mh+/hSbxJ
/uwC016sHYPiE7Moqc248QMDCFhU5JXtbb12I1oKOHhFOO9KLGIilwTNTYo6t80ET/pNte6SmSZG
l5LTW7rGdqJX2Rfm9I4rLhv/m13Loc9a4vycul5irAE/UwNGArK+lmeAyqzyepdzxPBZAxzdLErq
DsMS06ugiYDloMQOhHdEgxrVwZdHk7atBTEpIKTWt681lQmeognX5wr1bt/i7ByLRCApz1PnJg5u
SZQPqgW4Aj6X40JR/iLJPVtK1H3sTyWsH5AtxEmnQY8rVFk7ddw6wVU73BQq0uyomX3ISbPqfTmF
HqTJz8HmMO8U7PoKiJ/MqHBbdUPg7Ts0B8r93xA7FEbBenAScyEr2L2ltDIAVsdZVD1E+uVxE1br
fvwWJNeg6zRr6yuF2k18p+IooE/8JKiSDyBYZM21WmlPCrR3mipeHCTR8Sf8hhwe67JiOfEN6JBM
3NbnunLAfcrPYgdivDZ2x767Z43gfcBSL69hV53moQHKr34oGyNN9DJXVzsAjjWKlnNKdfOvBfap
T8Zxs2S4eXvXC7DzAjWHjhpkwuD5Y4M9oaLcxyoe1kWrw3zqo7TOXq4qyhut4oqqC1Xd7oSorZMu
H/myrRcpqsdiyY0LozxeCWaIkBFmxriVXgFqXborAUmioMYJBmoomwnPNiX/KonWTd/zjUUkugqL
cVTAbhCfeE9TlbL6/zh3823tGgcHyGAyOInManQHQGrnPiAMO9CicPXOMztvRZTOJsHY6j0wSNjo
/rlPwptP1+azkVQgktofCNvxuaVgjOAlr6ZibREu2oLzjGsOFKYJDYgiaBzAiRDtjYDAmeUevxke
rOaMT7lP4u2BlRHDR9U6Lplr312ZoQmIB3nStdB123QuMq36E5ZP6272iU0eh1ta6DXTgF0LC1Xj
M46eSk/D0j39K3dvKVa7lJa6rOCrk2NbB/i3xbkEOtYC1jYepLRr+7EEV5dph3JpG4oDgjuDGlB7
VbFN0rpRarNPM7pxHvx+11yul7OYEsvf/v0daRVD96fadW3CJ9IfL9ZTwf12PIzGsmoPdHezxCgx
lU9fmK1b0l8DtUgquYB96oqKXf6iEH+sRWQ1T23gC4KO9KRsS10SLBKTnqZwwIslphylccI3/l5g
47nL+IRYFNAq2/Rk6oCLbvq5n4OfFMUHKPFx1qINb0JXPvqF+9qdjFWPWDhUMV+93KDB5Cud7DAM
9hGBnOOQpHIK6NjrHgbDDl0TgN1gWwOVs32jZCU/M7zdJbfzmWQa2jRc/A4FpdqwjMFPDICxkbjn
WZtL8s/qzsecZ9de90yIOeJ5DSwG72sljZrq7LuZBGqubNXBs5XooJEvCCPIxxivfmLGvPaGJ29o
/Mw7ABBtwgahuKtQIsKPfbZW/3Pv18YDL7/OhWw9zZaqpoLute5Usk22r8KaFGhkW4KZFHuiuMEN
6KqpFXvA/mXmxFDuX3h7WnKV0Z3G7ONUnVBgK9DkVGBVu+D8y04g7Ox7Fz3/LBQA9JOV3hjnzS0S
pNwf7YxaObB/sgFt059wQ6rztDcJfln23o0YBMqIWj6rFlBLrVBEHjY0HkwRxEk43cygjMknyLzX
wgktJyZzzlrdU5aozR4umHpDeUXBB9PkeHtp/u3d9RYxk8zeOCPeqPthPhJiJTsRGZ1qTeubqIT9
6Q7YACAQve/fhiM8XVffR1y6xDH2vh40rbqCLWqoaplNxSHtj+V5MaJKAMaBf7Px/i406tv2wjqU
U9IYqVvkaFJPQHVGWwt66m5K83Zd/+isqfIbOXapWN4qazLnZrmoTr/S9Zixop1j2T5BYKH52Fbt
NXmv3QgL/Py3dXYnYMew7JPIuCYDXuX1LPsmx8hyuUysbRp1QA1+957jHMZGjNfd7FNbxB95pz5E
Wfrf2QZ32v7UgyRwv7MUWSnKHiVTbmIDuS7+x0PWrzIU1HXLfbvUBebeGKruJJWMNO/goQUggKq/
jGEohhnLDoBCxyCodhPZdYKaBEu+ZmSHbMEZJAAixVZ7ClDRK8RP1tBpnduHdpsGfGY5hzeXlO/P
5wCjKaLANb3an9/O6vW/CLO93nGWbHdX/vubyM7hvUlBL1QqbRIjEaiNcCIprVT5kP9Qowsm32xa
dAgangaOpiCKmMUig9Ab+xDj2NrDh8SpESEerjN+1frPWa1fmoP0Gr6lzgPYyGIaD3M781RjhjSV
x/piJgX4WL/E/zTdwD6vpgVMmMAPIuMhVsx1Cgzo8aVRepFTXvu/ylOaJSVCRIlzu09QQxSOriUl
ee3P8iyCn0+CxmSkgOU5UoCb4AHLQOvYmzk3Hdl9AzkBmNI+tUT6pbs7J8ar/eDEfwkSi+LF66ME
8GAx7o5EfhCRR25sfscHUcmu2dDDnsjAm71B2fSAgMMy8eWDVXTSoTUoxx9iiRu7kwUjdNn2tPT6
4eJSETxNF2Fj/wUt7afiKS1nZBOHOhRKw7OfQFtnnF+8hDnc8TFdDzGvgvLF+ph05HbP+NnUMIiw
OCzOh2sogrthEwZcTJJvcSzLYf54sNf0ytKHmrfNlnMJna1jzc3f2DuEXr6hosbNsa4oU7FR3eQa
hA2ujE9cqoX37l7R4pSk/c+mWGd71w3lBzLaAc2rmRnbRRdJmt9SBqZ/34n97wy8085CmNLJpLJU
U6q3F+Ia5D74SH24bPAgICEz7WVBreXWWguP6fL7GkAVQYLRUOW+6QGXdCV1uNFc7rYrianwfRf2
sDnaC9uaEAP37ETxKP7d0WjpSDQMHVFhHBq8Ob97tHoy8L0YFQDbYwa5lQXc2vFKo9FfjRe1p/FH
Z6Kk1xefsD7rRJHzfN/Ch6JIpxjcggxwbw4ip7Ul4c7I0wHl+6ZH7APC71+goJA7LALvS9wMfTSq
uGVX4Ymx1VqtiJh1A/VDsJGbThGFElkJcSsKCgAHlajWk8LrFXZcyZ0MXWlMubTGSsVLeIHSuKX0
kYIM07OUbvBJRMvkSYiktF516AWe6wMe2um9s10EKfGLPcsb1Ejr+OO5wS0HL3EIDykT68Nho8aL
xij8ggiTdbSqbrlv3iwchkjPYla3FFmvABJY0fWy1/ex7n3wT5ILMGx3Iz9AXBkFyn2BL0QKm/b1
wfzdS3E6qHAv5v9KdyGirsql4VVodkUBaXZgGm75MPeVy/UL3G3UK4tHe9izWE1KSw45IC84YYCf
yVKi2HVfFVDGNd68MvcqQi7Lv+qnt7Cd57Hs1vEne2UQIkpa8bBR8EN2nWGquzb46j2xy7itD82K
UFgrpbVXDDUPKLKY7bPEWgXNmpNWsFHY5S//VGwNk4UIdxMgcjajMTrX8Q5EooCEhK1MzvFNosPs
NdnQlgaLOWrMFYs5O6LTL+tNuH0384v5+35z8O1B4u43EiX8rJSCz69kLDaig5AoeRGrSZKe764t
PeGXxuWDmBKVZL6s9+QG6lkAr5UdJfOInti4Cqngvl9usnIMkHYOuqKgEWpDIwg188SwVbHnWqNe
YVrfTytwGo48DkWlyir+gKVsRqQYuoi2ACezjXilF9vPyjrnhRFGUaGH/URAAUfE4RM7J0NCev5a
VYUTpg5tyUdUiuU9EKFt2stPXN6rv+3H29/9L95/1VVrT4Jg6JF76ICZv0UGwce4egxF7CejeZcY
aY2/WJaJCZzDLRR6xZpsVqtJLqkGYUeYqtELLuDhjxlG7ZCUBpyxY3x7vTge2BDjB53NkUidJljw
kTvX+20plRB5TJ96rpoeWiHDFrZtnsNKfVwyh9kLsYOK4W63EmrCh3oQK0LCZikK2ORv3lcrrmee
K2E9UR210P7ysDZIsFF6ieBWxd+AYP82yCUqvasYU0zUST7K6iQGUDjHxjemJPRQwsqEKkifli4+
mK2xh4RXbqxYfz2crjEMZ2wvmGBM2FCwTh5DFSG4w3SOMKo/ojb3v9w94w5DWTW9qJ+Rj/sz79LM
n7wvmBvuRi7W0yIni79oPcEu5jrFWEOQYyotXVhTF4hz21xnOWC/sqtcxcs/FgZ7U8A8IzwF+C59
SGBreIPPiyDUKe0ScyaRcIlYw22MpEwAuIiNTRQSVdrJ/AxwZdfiTdMkwD+d47Tbrys4QqUYygkl
053rw16+aT9b7sHD+Yxb0PkcRHJ4t3Zn0lqbieHF/ynlQ/nhunEAeCdpdXjAB2bJgbRL0ukHVxzR
gxRqXKOtUjQL/gDeIiAf846InAGdv9RPVe3bnqNFIy8rlGixKerRk8+ANWrrC48uMp3Y3c6PK4rv
ow3QLrEDMsElq2qsJhHjmvk9sPrBUcbkDzQlaLw6l48wMDCrj4J2Y6GhdU8yZLZ4rgmFK+DB1yzQ
hxqVanOwsYBkqxJdo6cVt9piaKLkDf6TALhWEdIporY/lTzDfvVYU3+e9CuOiFXl9e2ecJcAtVc1
wsff+lI9/y+XZ6+wIThZFYtHXAqLoD5klVufWW/PJoLKW7r9A5rCJ2V423WoqtBXSlbqVMJJJg6Q
PLxPBrUJUyOQKrQpiSlTaf3jVSoWKxDVd7g2Pii9UZBqaWeJyYMTF0JftJGx80qrIPkPbKUnDqUQ
9SvmA+MZxlwE+akoBBTndvR5zHR7fNeTpXJ6w84xkDmgpL+Z2mdLw8tk5U6vwnqcrg5uaWH5jzI3
NXJuM2/ovoKKjzIolssFF5gNRwS1MLKu9Jp/UK8G0NgoEk2aDuW/5+iazBGOdJS56+jASSt/jlaJ
2de+ujedF7m1VJdkDHzLFMFh+hflTUVtmLsiiACUTRpEioG4ImIdUrq8f46imzqJFVrDpT38Z+V8
4MHpTBJ2JqyHt8RK7HACwf4NIJEbPHt9AC/9Zf8ETlt2nPFP8cH/Pqtdx1+AQh6wLGsYPXgk1ykz
9G2wnlNC2pv+cy1NHuzr10QivCRUbu+IbEbZmudyycnA3M4owORgGmjdkEL3v3G2hELUxEVb/J59
IYs9uEgd9VXN1W841PZK3XBLH3jFuiNpMqrAZcUJZgH1W6199beVt2ceLPEquUgso2dyhCif91U6
u7UJqo5zayeYbDJH7k8MGBULm3s3mNDkyDVNhxhyXZG4t44boIrE7pthBz4QkThMuBowcTNJLMmu
0dm0EGd3zLVQ0Jxj0jANrgaQIAtifivc7vsluEqRx0gCq6IBN/NEJEbPn75+/NUiywKTBm69r5m2
HYOWrtGKTNF4XvPTJbjnemd7gHTzAM/XXgD+DeeBJVHsMh5zUxm7w1tiDRu3EOFI6v6XHMXq7pLq
qnLnGjxKAQf+X3IpttnlkQIXKQMG2948E1irBLaJagkSgogD1U1GqQwyW1Uejy9L4aGToBnj9+rL
upMyTwb1PjR0iEcCcBgvSvSe99grJUAl3D8g66XpgP/A44ZTZ73fEe6dIlCyXhgqezrBDXC3mMzX
STbHWC1NKpbDezdQZa3D0idRotdmjI7fNMAa2E6K/+iohsa1+uCCOm9WZyAlv50vel7iG4UzrILH
RdS9RLs7Kuz6Lb79e4Sp5Ux+Hf02xc2nm3o0AN7c7/nSKXbzKHCuE7ZE0fMaqkSCh9S0F7ylNZ1s
VzvgK0MfOQvz5FHiocjLKtnjWhZ5yCum0A0TwAjEUJECWH1O5YLNZFJzjo9ZtNAKaW83N5/JQm1m
G2l23oFbFxIgjAx2+Q/UDG4IdGIfDtgOcOlRLs6lFBmWmPgxzHa6NVGy7pSi+Ego+Z+knP3cVI7f
sbKLfKtxMxzZFla14Wtl6OaWcDhryddy3agbCOgMm42rn1FyTFW4N9+WE6Da9+JzSFCPuCpU1vbu
WcDlyNifSRQzlWvNN6Nq8e9WgzuVt0O2ZRDhw1M8mnfjD/86ovfxmgO16zGD31j/Mt6qb3/yWvRP
RgsqJIzbwXNKVEOioX2jcHjO8Wu9PcPLdsiSP0Se+iY8kuk6SavEba0K3/gb2X8OKRB8iGUeSR+T
8/hHjJZ8+LvtrUkpG1WBHooUGXWqIN7UbeGHiREosnKjdEqqfoIlMu5VJ1PQNsigMdUr4Txbzxzy
Dpc6xZTyHUe/MIPjlFFxdRh5k8UYV6fGH/I4//C++zDGof3RiKVQDQ/THYgB3x35wxb/rdyfMF8+
HAWVhpKlXu5YppreusQjm6cIM03lX4FNQcnKT5X7y5WMC+EZxmn9I8AdnekeL0AwfVNzs7OL9xG2
sTN2PvXhmDZ9Yp9BfuXJOnuud/Ymvjkn3pjIDz9jO7DD8+xfkRVMJ7+blBC0eW3QD+IFM/noKrOp
tYjqB3KtqoLie6sf0aLWbNh42rZHasBUK3Bc7zt68RvGWTkg0oL6e70j+NhPl/Sv0+EW1GC1a0Ep
1xXTO+qLvdvyt5HyLIm6Ei4uoqG6NSjMRHXxG5uSpIZ+ooMMlQDOe7ocnDyrjd6xqAK2Rm9BRYO3
cCLa/eF1VSbWgxApEd8bCaXOC6BEiDFVmw97iUtR57nox6knOm/JVH+Ym944dt9rU9XcITuE8hRo
FP2K9j6k3PcxfAoFPRxC3TFP0ljHHif+WAA2RgGJL5AlUTn2Hu8BwJvTZjgwBym14NCSVtV+7z7U
yHBvVfeXqegjQ7fbmI/mm9KUVCc2AOP7AlwlMD/x6l6tx3DBzcW6uQGgfo9CERbBfQZbKDFa5ix0
8XRqnuix437Cdrw8TQD4hf0epmpr/s/pAsR3LosgHv2IB3JpEp+5sN2xDXFP/KoWDQewkF8Y+P4u
Ivg4KlmU9bm0Tz01jgExXRzwFXYd5jTMXynCL8/IBuDxrOJvVPD5kMTjTE8RXmrRFvfGIv+cqfTr
w6iD4E+fkJSWKJDyx3KqGSrHTRO/Qila4A29MTFgyZqQg55gyGfSwRefRokOxAttHctkpgLP6LS9
7hmOKGmu1NdOpEFzLf7+getPtWNGr8pPcB7t+ukQFN2zzp0rgChBgmElCP1foWCNwqILxob7Jh1e
OBhRhfvdYy/YXN2pDzG4bGfSfRCRUrY/2JGEV0iOfA2Qu3Jf8igp5YLZTdnyq42n9AgxErGWZWsv
uAGideotQtxc57kbef0s2vTANYh8km3gxd8lQ5piLF7vCzh+hbJ+Y77UBlTyZCQ1AXezPVuFFH1f
95B7w9FF9Tb4K4vI/ioBtEBaqslmp6kzfUj8wPPFR2zXDYrdG2Dr+7DdCl5tEs73gwq/aU6Sv5z2
9YmxNRgdytZ7zzCGcsZPaZd2bW778Hg/k9bb+8zXikofFqkEm6tKnKbnrXLMlwE/C99mrhOWHvp4
3uZ5eY2OVJf7Yi5/AAsbw4di2qVuQfUYl8NF4HyHZgyoZJGN+IDKaesVLTdt3vWhmo1fgJHn5YIZ
DJvOw2SU/5MtGWWmG9rZwhRVObQ0kYdWLMVYeU6h3KOdpc5M19L9/AU6aJX+RWDGsMGHwnMX2rYT
ShMT5xeYA1a+O1vyaZnEvq9AIHcMQNwPkkBNCx5W5wZKRGU2nTnnqgHHqNRG3TavzWy6Tgurm7mz
qsN15tVH8Clh8B0+PlKQpSSsjJVYo28rBMQEqrKaau35184GZ8vJouOgCD5s8wQnwMeSchaCnUwA
sGWUoC0LxSJ4NS90FJSQaa3GKZSKfVvQ20zeJqlumH+r68l9FU3wx2aBMt/fwPHrNYfVkN/EI0oz
/ru1Bezr+/L8zMbHJe3NqzdFc1LfRuOjgqScV5e3vOo8Lp84z4y0EeQVjCLya9WyQQ0j7ByXZ89o
G9eiYhFSo+Y+c/BscUfgNFG4a0d957TvkwZvvZNNyn4fkZrzlq9LEsmPmrNlpfLGGRyX413tGq/m
fg4hOo+0coK5CYn/CiErNNohHe/8DN6ss19bZwCFG+6AhVw9Vm7tWWF9Vhwl++OgLKxV7KwyW9RH
pmsWVm9INru1LMGlJOyKYe54PLmuSIXLOXyTEahsZORRj5Ms23hfjv/4n9snCTCsVeizEtZM4lP1
+lk5wX132fDtmtubvMiNL3WuaP6oCxAAmohvIoMo2xiIJYz04lq27kYNgDOwXW8BJUxBFBGPuzSv
AEabSgUc+8fEOCoMXwHwLt+16m5DOJS3YY5MdnwSSagCxfUohBqy3vaXKQzB3Dna7BhSJVAQXCvS
ZebjtNOfgy06P7JhGW4RSoHlrXgRr87Bh6GSiTdvkC9Y945uM/rrpMAqZYgUYddDc8/oepIslTeE
FZ9kCDetbZ0EIb0bQ6dwlFpiV98VcGEDjj08yuMQQ3GW/fk3tJT5S+KHM1KjLNbk2GoPTZpkXhI6
8vEvGs/NOJQqkss3dGuiIBwMI1Iq1HOXRoGDcfQLHYgJ60eyeNAwGopASa/xxC2wfjJjUMVW1otJ
IOTaimiYDk0xG8QzjtjQs0NaiOvujwayFBcxL7oZ+SZ9eUwvTPZ7ZWTGdJNzfoUtJ+NOXxoHghfA
hyvmhlzkcLl+zLf5OQyYhCApYZU8sVRSJqlZsN/6qbyQUZ5MgInmI5FW0MHYnyG1J5j2a776wsPz
007u5mLpYRreG+wSTKvihUM1fEvdPkCDpi5XA/F1DuSBYcfvb/14l4gJiIfZBSU3NhcIOEmwSCsl
4Dhucf0Mw6TUeaJ4Kr6nuHBD+MXdJKwWSvg5g1+LdoYTUvIWJ7vFVaap5CG8cEqsofQ3ns77DIHe
ndQWZ1qQvXSt/7axMxNwGGPp+rz8mjxhpQtPMEJaOJ+8u+iGcgMiSUlOf+tT0p1g/ttc9+tG3910
l9vjoCr52m2I5LIEcOPphZGSwoxtrHw4VbXZmIzFynveuQbZnWvwPr5RSf04qesSsFDrNC+4YUMF
8wfRPG6XjtXzaQE7Ae6hkCSaH7sXDEOwUe4P0xh2KnjTHZdUWTDhMKqWRV6ShoOZpMj5ecA9U7hX
KLDEZg67g2D2rtHtGdhULc11u1nghGtM1dSRoZa+WAFbwC4Xf/uxkCblxs55WpNxRvep2qaaGhKN
Bnwf0ajHNKQ02Wkw1CepRex/1myStnFEK88oYTaKOt+iSvc/8cLoAgUQg22+UtTBQ9FUNWsYY2D1
8pnOXCFhSvMbh+m1MmwcSK1N9SHJJO6XsRpHTf3cmX+81/5dgq1bSZ9Ongat7RNYzG8tjOGBL/Fl
1othTYXL5tEdzYfn8OdbQpXeNqxnQ8NBHqJo9WzntGknxtjdc+zgGeUtSFPHs2qR6w/5bXYvWLeX
/Yy49spKTpctHopaVrfnJlaEkj62xJXlE75HRKtdkZrEN8kypXnYkJw6DWmc/zsqaFruISuRmL+e
wMerYlX0S1I7fr+JMYEYrvbl0/T7ona+6M7boqvJ7yJkpa3QaiupD5BnAdmkg+UVTydD+NH1I2Hn
QJNziBa5SZIqgXo9Dyuw1qXyQMaUpFhsQ3ZRJLS2GDjxd8Z6S1snoKTajnUtgSz6XUHUIdJ0C0XH
Ks8N8YMlbXuyvLfcfiUDspm/7s+qjB4qVUnvPHAy7Sm8WR0jW4C7K5jnZk6Cj6YjkBTClf1GNvGT
C0sZf6VTNJ2D4E8lZ0bgxISkZiUmVP/Ygm5boo/QAkeNd8WGT/sIb14KzH9wKzlFezrTeu98t8Ae
ZpQwVgJAcc3tAABD8o/+dHMSW4R25yXOCO4VQ6Pu2zg23K5Nctij5SFbfu4xJnQs2yqmAr1xy2K4
FMDH8W7ACW9G6drBTtEVKKwYLd4z6mv3Xcydb1d+X4BsmLs21G7m+OUbA+oBGiDAGXIKnbwWf35e
dgOnnXR62OlChFgU5hjH0/wB6R+tTGau3IdXLVW1HxDmPNT13L+UKhEtOjmf5HozJ6KHGYF9EYA4
TPaRTxKMdisfzX21KlJSKq+x/O/ijun9SmaisoRpY1V7q5HaDCFQZh/f3v2IxtJNPSIAX42qET0O
vTQWYIWpr2WnPUf8IIvI8Fb+xb/sAs7rS3tWp1VbSB++DXoA3y+68cnBA1D43sWjOb8L22VlFCdz
OfTaWUizn7h29CiMzZcskU1aj6/9A33QzvaA9ww+Do5vipbBjxqtGFI0Swtn0HOygXOkjGMc62Hs
1mnkqV6HrAAi23DTIYU9sV4IXHvu3a6V5ecvi9uRyjdxNG0jV64+KyqG/3mQl//aF7viEBccGSeB
Aerx9hvz6o4EYr8TRM6Tmkp5Jl3Fq6TXYmdk3UPlnhhZAGvBST8wPL/+Hc7OONMO8dssclOaqQuE
kc0WtFOtnLik4HtNhcApEOA1f4bQPS0GcnNMMiaEDadVHJHaVhuW+yknI+02XrrGRa6cejwAEtOq
beytpm7oADLlYMQh3lx1TdZJ1MnBaajKBo5dhc+9JfUD6TdZPO2JCwArrNehPR4bXxu5mEkU6w31
WY0pJHQjmV27yVmdqQy4uuReobYeALX0Acve83Th2xcO5CqYsHgBaX9HYMvNCSjmW/1wQb+Po4T7
A/QcQ7c0u+r02dCsGp9n03e47Uw3subdd2B7kCLwSPrpx7InDRHwITGyWNWczx+iK1n99CNeMf2K
VcmVa6vC32yTD22zaJ4elTCXbi+czlquCi2OTHgIc9o3wVWwzZPZ19Aboo76YQYY91VstzV+xwOP
Q6lpdYnXtQnNk4Ed8FVYGiV8PMS18YtonEi7ZTB7oSRYpMst5H+NjMt5gUrOQZHL4IGpJcjGvazF
Aq92o05rbemloH0YkNKNeuaMIE0p2dZCIAAWRqgdriKB9e0lfeO4UT4je9AYDR6hSUd0CYz5Xrxy
fONUaj2RJLb7tWvOMK/hLZ+ZFXwiV28FPTFgkIjfCs9hyc5GzEyEyYO5mkMEqrVKOEdYPi8nmS9s
p+5qBjAuHWYnpxG9mqEfeC0Ion8VC7Jgo1xneZlJhnhlKauyl+kpsmxZOcvRPwh3E9cTw4ZjNmrx
Jb8RoDybScLs2FK/XTG1zII6pkLxTvNj5A6zIth32NzNwYGK8rKI2tSLw7f6dWLqrCLe2yKcZYN3
Mc2T4oL3iRsGBbrMFwUQBmPMciNJHMvP8XlrKIh3LgjVATiN5C+cxVsZ2dVHyT4aUlZknP4WHdWQ
dqkqZlDF1HHjzppf5N4IH6bWCntW57TpmHd2ZNB4+YQo5uJajhOpUj2ehm35g7Ni3yviTYkw9obO
WjtMa5crlZ9x3nz5jIPzEYrEhxUL/W2Om4J5jdLfY5kxYxLKanMWuV7yw7nlgoNKzAXmRI65aAGz
jKyxU1ap7NWJKPQNQcux/KPj+SdCt9HkdFXolGGWAH6TkqajNSrz+yCELiZF3XADvRThZLjZ6Z9R
IPxZ6DbAyoFGj2f7kPkH5ey5n6nQeJOWo+XAkcDt8Bn9Scg+BhZv43CLxW0/F0NZrRwGBsg2btsc
ml85LVq5Bc+OmAYMxG3uoqvY+pMZ3afc19MbmhZx0LPnEEyr+NztkxxqtanwzwDi/uB81hiwTJcm
piqON6e9XueZ0ntjFTz+IYeD7bKkX8/UZ84SDcJ7Erlt6oA4tONfWMK0JxAWmRj7RcAEmriG8924
mVu4Dx33ckhqtlUErAJxEVpx6Zoj2XCHnMJwqOH+RbHmwtlIOX1yULThe2znlcmop73dHW1+6Gh5
u7V2ZA0e78Yn8+ObD0dTeA0+MBtpCA7Vc5xK6h01Sggjx2ryXTuc/p/D7d6XQuCnjq0paIAHXgaE
9M55YrVKWx0nW1fy9olnSEdUORSkC0MCqcV6SPDyuGnBW4F3Jb4R6gGiMLm/RJxTsNEqtjYjLgD1
YGSI/Pg1uGS083H1vBNA5J2d9u0D5GWROZyEBfoVzugBqK2gshoCBosR2TZW+9FJirMwhyy5w1xY
PS81iFZn1SB+SJ6zrdT0ixJxSX0VuCsSSumZfhsq1bPEnI1xVaYg0VtutGgrItMMbTewGKMMiwcF
Abkmy+Ck4OzFZiQQ/lJB1MfyYimaJdKwzpBDRpkytwKB6apvX/mZzisv4SKAdU9/OqdDOa44dmza
2EWxTIDg1NUGE+QCFkYnFyC37CqkJLJw5r6TDmUz5YsVOmUPU3B6A/NqCVN3HsoQaYF2e3wThLdQ
birfBYxNzSvIObUGmvl6l5dfg7NXLTNY92yrBkHxDAase92SceSlrNRI/cGqFGS8EtCJASVE0omG
fKtCWJpj9PDsQrw0qhi7iCU5GXpha50lNJmrPvLXBh7KzY4xwkm6zpOyE7yhhU+U6405EB3qJYtQ
ysnQbAnTOg/esPwkcBJBefWlBxTZCrr0AwACQMvxGo40pVVPORRW9l+7EgzEI/QLMXPZSXp91d9L
MBOcsJqEDfcpvNe1jJtrlKZMLWGy9ItFCzX8jE7mo8/9isOWS9mAsbIUV+XuW6otKKh7tjbCPHvu
3yO4i6X9O37l2qEFb3DC9mjbft1ydbOegTjWOAn2wxqNxO2kly2HhucqwYQDxowvuUm487mCMf5Q
l/yb8xkBrvTcfKyUktUyWZF0ZTfWtI7xrb80QphfCTph7SmFQM2wj6QlhWonK7je5GNiXSggeGkg
gfFkyoJ4q4mdsCtAsyiiZTc8O8M/04O1e7YbgdUZGUc5YpK5sSWS97C8Q8KhwP0GSSLlygImXti+
mTDC9JH4FuHLqiHr4KhMjg/QVLIRH9M++HrNtS9WPOKdxMgeLbbbQgBs7zKaFZxr+n9qoAzSdqsA
nKvz+1Y0cuRpg+xCOAo8tkuGJsuS4XgAJMywctw8DdUD52GeDQmrukwwHXFCAHjGHhOwioOLRugC
aCZNUSHcBiZofEID0TZVYwFBojAux4h2Nf2l642PfhqvhF7ErJrsig5ASUuXZxuBldlyZECpLofh
QkTTgqCuMajNJ2NAVSYp/6J4Kk3XfG87chQ4RpFlJaIGM0mmtteOjrk8nz8RJ/8N4RTG5uGMywE1
20nJDoeHps6F7UM7XLrB6EHLMHPGiZkfbzjKUq/t8+WheUDjjYKUitufvIUQy7l1F2r61ILrImfa
VKuET6FyEQe6lPrbe/x15QSR46ZX50aMZifVPUUyVbkre1P6XZLIA65TDYj+mhG3x2it1LCs1ni8
q1MSXp1eS9HaYyjqDqmFpEDuEpzIiNdB8ufsLLMk2nk5MoULJUfsFQkM04gSfL5J4lidoCqnfeXJ
Ddzwg3pWS7eY6oVeouOPgDvtuXvLOiCKx5xaMLOtR9Kay6E+QcejmyYCULNerWMVHScaFtMaUanf
yrg48lrZ4+i59h87JentACHc4WSRV+M6Iagd11Juc973+VOy15LFMI74R/Lhv2GHcoWYYn9YQ5qU
i8UbAiMXj3wF0XCfmAbeFCaaQngPtKuMV0byAxR0f4uWKc++7ZqY9qdq3fbg51fvwRi8Dyy3DO1g
dIZ4Gmww1JrJJJ7AF84oRi4j3kClRNQKvujXUo8zZC2n4OtH6hrQEGkqMkq2jhVVbBWgootY1Ks7
xy2eTCZfVkMubhg+eM3ZPSsL6xk1FscSz5UpiEEuSeI2lNPZV0twzAOBJGJxER35oBM8bOPiYkUb
0RDCYNaZkyryJBiDPwF3IB+nMFRJo9sFy9lUoQmdder6Ci/Xq8gSultZBfbUcF1dk+xT70/f9QwN
JPaDoe5ZDlvy7qml+LdqGUdcC93OjBgLANgwZRSLcLOmuSk+/II8+O9xpLPPJETsXuZMvnDduxBY
xPqdPOj/bYAO+HvIjcMU0bTW5yKEdWdwj5FG//PXeS5k4qAjVhNCMrpmPD1qKZkWiq9Rdm7FnpJf
zj/HkUQaOHAJ9ykkxDnoU1a1vEy2PByVCRsaxRKUV4SIXdfOqsw7+wZCRHoIotO/duxs6kBleRNj
Mw8WnnQPyNvqWI17nCxEcz3GH4hwyumr09kpQT+VBB/qYLzhBO1D0WpgC9joTOxRmwAnMcDaxmpm
XsuqeD2lArGOK8de2htzLaeZpSmRixiqumh+eS13Xs5eswsOeyhdZZsChJsOPypdhfF9EREBsbSl
u+MGWvmcmFtjsgig0TO1jYIjhU/Lo/6d+v5E0tTPzajoPBMHjHxwsI9b89vnABWuhnWYL7qm/oiV
aoIBUJezQC2w9khRaE5o3tgPUgmaIfbrzfxsCZ0XbgCRvjR34FYDaxdIvaY53rn4NubrU3R0ceUs
vK29461exNRgm8hGstKx3BUy4WOTosy5ZK7X3wpMkSSkdu6KyIao4n8AG1mKtIbep2F4iEVxV5yA
cq0hzgkp2RZJdSqCfTpGvYenS+ImWkdS2kccr5Bn+nNsa6GCNGklBoSHavq5pUGnklVKWFjsItNz
CzQYbA5NIlanRQ/yrrreuTeFr90MlDMGkTCeZk3cAYze4clhfx1ypccBDEZdIO2EuTohHnqWyvkK
WxmctElqK0bIxnnzrgz063/ycMPjKN1X3jn9GqU9+RRgOrc842pmsZhdI1KkHX4MxBdQ0JCcSa0p
zaJziFVyNyRO2G9PhMqqQmUCjXViYQRxY5UKDZIhe87apXniwyB5LGgzOSfVqHGQXyt1ibvQbeVM
uv9qcH1p0N+cvUCm7CKC2L6h6vYofBsq1Q55ioKBW9LQLvsMARV0nbqnzmukRq364v17WHzgPVob
vbm18Ms+ZCxNe7jDqfilKJ3r9LjeCTK3wf64BIdOMZVcxDWIRoU1pAf9GQnK9ah7qmxVmuGWcb3O
RSFWfNCVXDf3k18BILjOvy95bS7rFM6X/d0VBikXURlay+xf5BTE/qDb9DVKcMEO+9wMW4UxBZem
tt5MnTbBnAY/9c3NZR60Iljw2IS8DKHovoT6gsTj90mL4OhlLVdw1kQ084vlvsHJ74VBh5HEMIL0
r2NE5KtNhS3MTXf+AxgMT/dKJY5+iAfBszc07hsDlArbEJjAICxyxuUgxpnmROR1vN5c2iVdY2/2
gsEbDvFfJb210tSIbua/p+Td13s070i/f1I/Z0j4gKHY1ZZ8lhhMDyQQzdcrYATwR8F7tYH2QW6l
4ztSlH+KqjNAtvP5vGrZHBk9X9WhVNa0vP2HjOoA60LV9Xn1zIl2jvf9ScNF1cvDL+IaJugQ6a35
gquQAe245qMdgNHgyKO+9ym0ZMH9sp5mACJzml60WNxZ+XXzHa+OGsjAOJXzkz/78Mkrph0E+1I2
oPcEac8Hb+Fe8swWs52bKaFQJ+6cB4+GVMuejvCgVfIGClVIVFtmUwhT6c+p5UDXxP+fPnMde8RA
jv6g73vSOF+jDgplNVVbipoVaOgab3FGqzC5sOs3gB65paAuvRVxkd8FNl1kRxET2uM3tqVqKplf
9oV9OvJG48sX0eYvNOOVsBBA67nh8HY8lkPaWSOFLGcGArfOVbsRVgOTB84iA0SFN0e5iqIwUL5V
ohZoj3gPLwFYfokv+snNaVyoKxb7qC/1suABJYPiqwKIbRn6MHxXunsADnLW0JA10zmNLKwZ9tqw
ZnG5G5o/en1cYI7UxLcnpRSbbDiJ/LNEZqN/XTkXPL+RU4c5eGUuFJieOhzmMNrJpvtNasjd2Suz
kQ52z+Kk7RRbUjnqJofcdCuFihobwxVn/uKArgCpMnLcMhzgPNQ1+wLWJPtEUo5WQjTSYVVlO3Zh
NPXOA5Ek7t04VuImfdBY2HcNClurl8Ui5s+bjM/iSmmFz3AwPYevFk4pAaSWUaXVArLeONqlAh38
O1fkUO4RCaYdRQNS+6EPmc5fF+DiTAcPhfbDS2P1/LOwf9X4Csst7sd738EboDuT9ryu73Oz39Vg
qENlLaBfoTawRywou/FkmFuPW6wSZ4rc50oe0h4UJPNlYRuxkzgBqe7tOp3gK8deWsDH2w1sAv0f
X4Rjp+w62SYDSo3sJNVAI12xQhU+jZsMEhCO1xfTsD/cK7IvwZFObCVvT6DGoqU9w9DX0DsXaeWx
Nwzbv3j3Yi2UOIfvJVTQYa4FxsnLZxAFY/mQkjBGE1HQbM0QfqaxI005BSD9/72H0ONzCF5qFj2a
W+P4P0KjDRAuvsik3sYHhry6Q1j5l2adnIWG75JPWZP52VbvxwBIW0aAbwq1yJm0dI/4t2hF1jrZ
uHsrA457hYxEzBQwmYNYhpNa08fzTH8/tg74NDsrTfNbooGmBJbTmBCym+AEK+4OeFfCtcs8I85B
Nrj/FsGyyRracDYSDH4bP0EClMY/VqMdGahijRrgYgHPfzTSahfaX0T3PyfKcu457XKwHNCWb2D4
ufE0uBlW5gHH2oVLB6svnnGn6yfpDUz1IcCPNAsc2i89R8Btmk52os+ct513672JBYOtvlhRaicM
sH9RGhDHYNiG4WuHYdePn2xHQAskm8jkwzbY+XgFIcGNUZMwx7xOmgMTC1S/NI5ycuso7WJalA57
fNpYuk9TPreXcD2EnyPTNt/VBRSnWuTptFsoBgyUPlVr68MYwxOpntT7NoSmws4pjgsRd6JQHGsw
wVOI0UeRTuql52laB64MO1qT9GYbrINoON26lsXEEQ/XJaRNEzq4mdnGI8wT3hX5HDdFUcaye20c
RGK3BEeaTKZiNC2ha48/NXz591NfGWZAB7ZZg+9in5s9eGAWzKHXikJnaUMWOEVKfkJV8N85Yun6
y6hwFxu8d3Ud8o/RAUJFNsMbi7j2tyfSGO6j63g8zIQOkSNYuNPWn9KIZLWiGwHLwyCaCB2GI/ye
O6c0cgijXhQzNaNirNyQdFvsfq15YdgljWHFuY/gurKQty2h6MDnkG9+k4wD0rtBfTSSKn1yL8IZ
nG/Z9/ySU2UGQ2ugloD6/6D1XfAxiGXQ2HTG6gKhx4haqKWzTvEvG+K/4JvNrkv7v2/0TucBMOa5
NjxykhhW6yxaEf5g/ZJFq+oWnzqKSQ98EXbB37NhPuStX7OqPUMqV66SdmU1EHNYuPjC1jESZhSL
VamNkfUmy4wJVUD8grGD3xk915WaPcFFDuSYmm3BR5KSMD7twM08fdeIJaMLXN4QWignNtPmHouZ
6j1bOzSiWvBzRB3PLlNf9VvWp6ELmjf3xDeW3C1oWW/i84pnuhUs9OPRpdupSEkrlRoJVEE5vB/A
5zJkPUK7+asf48CqJSIlMwt5gEt91ouFGnG4QnusOd1pynQOFlr80fQXWKVbkykVTa1qOBI3tehp
rYYqkKVO6xLrZ+mo5F88fKY2js/ae4v/J1QIRTRSr6y5R6rJW9+7D+/lRvGvyN0A4CyU51RHON/k
7tIW2qJFS71VFJ7zMPqGMTzhnexPpOIRLQRfUpzj1FBHHZKiIMXzbKyorqE/l79c5jDnUGb+ouyl
24oHQlOEDP34Kr1ob6EkIXszt+xHt+S1rZRBB5g6a0zX7A/2yNzBdCupGq7stVwjR+XmIEeOujCc
ocnlM+Hg9yS+MustoZPtmCg1Du9/yJc5FTSGEF/vrqIhoNFrNC+BJ6RiPNDg+Kwc5TtlZFaDYG38
Uvzje3vugCQb7kHzpsZOSmqrSuowUFbHp3+b0ZgnE05s6KoFNGw3UENCxeqjORtG0Rbo5CnRQaLe
Q4PvArfIM9rR5hz64YFHz2KfJJtSIt1LJksCg6NOueDES0xdK2YsPh0pP2IXXEVB24E+ySzCfv0k
fj/T1Kj97Bu1w5O1NSmfAD7v2e61akdhKsiPEK/gHVj1k19zCDAvC7vqhtAbZXmuao9DPh2s6j5h
itgKcl2ghzki/5EevbYGrMM5ym3kAfvTN440MENlqYePmR9QvXlfA9RNhq1kLbMqUxHfRPpzcWvG
HjlYaTTnAy0vUlTqyTJzCqvGjlJtZmMlLuwwC0zdmOahjZTP6yIkQnwCRrVrHi48MqcZhK6RRCZd
NJi+xO0kEXxzHb/2425DrU65KaCLshRNosb4aBfc6H9ke9gA/jtzupUNWqiuN5Key6EGS+4et/Ji
7RR+cc1SdBHJuFoC8t3PMv06YF/WZBW3HVO4toFfBNOYJ8301YWRRqtzWZvAG45v9WAI0+kT86N5
LlNOCh+JwO2b605rF8iQgeXe778Z4reNH1iLTS5nX0zAGoOXt+AH/k51y/TTJ4S0YCk7zFdp4E+p
mqWK/e+574mLi9QN6bB7PRnEIMmzpLL5mNUICsKZKMFS70ZWF2mshxq+7cQdkTXK8j5hqCGEFCnA
qvfRJw1MhFs9FyFQ+37GFyWMzldjU6rpi96SLGb5n+SBEMk5P1exhnqeBIIHGvXIpeR3sbpfwXvU
WRJ/Rgk39w7b8rwMOlOqFqYw/MhV4IQB4ipbeX2CF1v5poFSt6J9VRrk02e+RdB3PAtqnuSgkBN9
dwPyMI9nq5lfT+sRxUNPRL57lsgTm0cwp7DEPSdLhwjEglPAv9KYYnLRTbjmI/LRqAvWjWC5eEok
rSbHiR3+SkT98kENW2o0IdWz300bpQ9jqFBMpYVSSWgOlHukNxj+qh0XvyemHaE7GwMXV8Hdt27P
uYx7Hnm/t73wSJ5ITbrh9n8EW5nHVGvqB0br66+yeJbwDV5qHuEyunquTzykfTqVi3Ch5V6qWUcc
n7GeukftCPY71kSiJC6MacvU01upyc57h12iQp6ob0qKWa18ntXkeFaPfEIpp9rkpm7jdLqxkjq9
K3KvNY9GOareRhZlkq4IkEtS4+dkzL7MLIQUfqTATcjU57zwNAPj+3Qql1jIswH/c1IFqRHfit3g
91c1b2ma8qdmgov6lun6WpDyA5YBhmVBZO0Fd9GOcwjanRk6bj8v/InE9Mb+cE78PHHI2V1/kTVk
SlfcJuHdC2HTPYA4NjRI6x/FGWu/gIm1N4HIuTFakFdEuUBE2d8g1mvIDimZ8J9dS1asJxFnQHvt
atL3q8h8AalIH71grELzeAHffuCEZOF03BfTUSL49wzdRG13lzyOTYMa1SFW9ZKG1vYjxC0h/rUs
RGciY/hSe/EpLNL6hGI6SWksq3OI8yvES/ye1e+aZnWUTX85JCPpDsC2Aa+fBgRMqUpBhxZYeJEd
YJj2z9G/10TMhNmFOhCSnSDsEmc9P+yh1VP8g41mUU6thsGMQn2DPbPhxaIiNqZw/NIGH3lm9APj
9kkOuB3XRhmSQrgftp0NTAaGJey/bU3mnaQCIKIsZWVx9np03VWdIC9IVBVQmkzkjNwpncB6EDiU
U3g6igs8ZhuwiIksFEXxy5UZk2hIn2ugHH9dE9syfRfj65XCgqnh7JHRarv53AJ1Nhe4Qhp/FXvJ
/uYUFqAQ1oVrChCXfFiJp9wnOGc3g/fr0xH/Zo+CZTvMoo8kiTw2/P7ERTqCG3PN7pSNq3hNc2Xp
2OqIi4Ckt++/0xnP+zg4/A7QAXsvUrPFqVc744Q+vtzBH5UvfoqifHqX+ED/2qRxrQ4szBwRYygm
4NFYIsHzKrVp+CVR9AnozynjHbDBDk/Av6QT5mNT+Fx6MhcAu+v4yWxNtkuODdmts5Z49fj+Ib+O
I5pvhJMWqlykZNn84YX4eSK2ARRj9uOHJBM1/cadzfrMItCgMniI/Wbl91doKwNxoaBIy/oiTHdj
lds6z6Kcdj4uBMtBk2B6q6hHuyfaT9vXQ1+q1usiJlViw8JnR8nRDRYuRXgy0iHCTSDNtRBn2NO1
vXmeOYRno5dYMTGIWlVwlPLgKhyDhgUkS1fgGUjpyixnZlzgztez+W/RNrzv8iaNukL/MdSjiOUB
GETQJgWhiql/jVFObjKRtdxrdQteRimrS9KFQum29lu/Cb8rxanx5RhXO7N/qvCueI1oCCuhzRp9
6/z2g/3PYVBd48cZuuiosTh4KdSoQx5HP63mluoXYa2Q7MBao8JNLCcB0u+4G5gP31C0ks+8cU+8
NsZ+Zfl5c8SUP2xJa8Dy6hYeYliZQ+HKx3BSB3o0gjnZSdz1dQTlLwP2fa6ytJWdmXr9APsiAXnA
71WYVPqYpGF+/BPJ1P89IAFdMDKiHTdovd8lBkZ/Sww4RN+bpnXrn1AzmuG9qVJmrczmf1KLhQqI
9AyzzLb4ciQwQQTqQCHcnY5OD8hBLF8+WcxAoGHPr+zLBL4Gi6RAhvUbjNsl3K2P2g2wQzqEQUvF
vRdAF5IAhe+RmNpwTVQDOUdyNES45K+TG41O1bSMPDgWy8QZGl/4fe7wM3U3Auby/KiKyEA3hgVg
krUiY1X9WA0fKFbaE5qSvHRxZpIPWz53/V04bIapjU4wtRtGGjQPkOMmSVFY+sMVBvIcU24JpZiV
HZ5IwCLanjr/QxAAJ7dhPFisttptv571pIhBpHhAhMyEnnE4aamaNYNknFrGP0+1fAWOo3fn/R1h
XPED69/WxUsr9J56QbcSO7Jhq2hgc6mIt1V4ka7lbJ2Cixu2OogGosvVi99lyStDmYyb4FAu/Sjy
ZxrvJ3czx31CSyU8ar1c1vrcZBEKo5vQe9stBnieljb33yI/230XAfQRSGwqCvBdi167QuGumW17
SuxQ95dWVsn5vt+g2HSENSeO86Qo2HhfiGEu3P5ixqgWvq/DIBdZmAfhOJ3hLYJfoZKLx9uwWIUR
gqW5HDBecdiGAzCnSbOlY0yyOM+7QeVCwxNfQTUd4nwt0Xwa2rTgpeIgm53bGEBhOl6Tgdrt45pv
FY3mQ1mvOymgP28/TnLX7l2B5jGM2F7Y8W22o31OwtUMyVK6pVbVd0EQKbFQrD5vDC1vJpmvK5q3
vkFZdUcWJphy4VX6W6Jq9M48oMRgCCyxGPh/akBN1MXMPCvckI5NwNEbGTM7g9ITFK1WC3ygVbJS
ERGtcIMf0g6SgjOkdLP++khR0YJM3rF9TrSTJqAekJ2uorPvdks0XzncodAsVvFdcx0OdupW1i8k
cRhMuff0wPm9V2o8WFSzZmeQN0LUv1WF48fcnp7vsZMKE6PhEJEhyqfdGZM8h4Tlctd00OEdDhE3
lGu/eIcS22j9SQmx9DdEXnOKEC5IlbMQTOPK5Z0UqskFWH3hxD9nY6iVYu1XfrlLuu7Ro5Jc+95q
YVnzrgSAIMTDQk9bef2wOsQWaPkpFupBHuDXFSpFvxnznlL6qkaEG78t1/gvZ6REq7pev/VW0CF5
P3pDY2Sc7gLuYMw+n+N8L8w9iC49unR4rM5mr/2ctVKUnNLpYfWW9jcl28qPL557WGN7D4LWcGV2
FEQ4x0aS0/lMSH9S3f4gDfm+BUmzoq13iiVaCwiSpo1NzMwQZNA3Ho9UmkBuKSYz/uIxYempRa+f
hsmnPZ46N9lqbzrbh6PefW9FYYyACGiIq7Vw2w8HSniOCRek4W+Vw7e6iQjJteYKdNauQ0AyqHpc
HAP0nsmC0+QaGE7KgAHHtwXOoxjKN3nPK9aBYcUk2OYLIodX03k6U60JYmVw318Xnn4q2cXWN3SB
x9hqyTIkP1+JsgXXM3SS8MMx5s23nHuXOPNL70xNSQ6FkPk2lMwd8qIGuo9aeNtgHbbrQ9+xAyLe
4ZiPOjWLlC6DW0IAc64Vhs4S0Kb/svcKVr0jPHJBk2SDHcUiTajJEoWjs820wBK6Ry7mGmSF3e8Z
5epVqVXE6GHLqyhb3Y34wxcaScjLeGHZVupKE1ruyiXJUAo+rjCqKHVLyJRVPfZHEcY3EHleXtR6
1//VS+o5WZadD54VFaOzunWCXHp8OkSmlZv6OVDMpjrq6oWeFgL04Cq1NGlH1rUGRiY6OgJk39zJ
zJuOsHMMnPpWZ9sn8EIRgUSh7bcaZBNk4KpeP4nJrKQSbQiqQHIJM3/39kTiGQ52+X0t4vNJPBCT
yzZkc++T+rAWaRbAtkAjmFVW0pIsLsvyzJjmxSTe3cXwgKmc/KKw7YSq/t3SROYaCRfJwo8Hf6oz
hDPQaNgmLVTE4bRFJopb5NPMuJDW8trP01xe4KwhvtMiHbPb5azr/RbYTB+5kMA68ZoR2Z4B4XsD
+tDyKZblJcw9ATh4r9d8WhunKM5JlUbP3scuqEhXGvWP55SYjdyJKIE7TqnERCyJpyVfEUOFHI0V
m22XUXP5095OQdL1R+3z5y9i97Go1FJ6L7rzJBpOt0XMZlcKWu6z6x6YXzE7WQ8iDOHokgVspzJ6
m7HNrTUlN8AiZbRAjKPUaKRBkybWhdBa/sDe4hwoRv+Fjtwg/hDmnaNJmFs/ILatSMvNipV+vh7r
jkdPBGrGqnFQ+WaKBQVUH7q88r5Xcm7zLgac9v7QjUf4x+4Yl/yHx7TZerU2mh+iHEwKBuNEw7+E
XWzXiOzS6ogDhd1emtBYllTzWT8WuT4DC5jYHMMr0O1am27uWwe9PSDQJE0svecoBF+p2u4IPL8C
59swtX+WfgQpPfGqtGvV0b2Vd1AKCSYAftXvkTTNAxNNOG+cWCiFiqJ/aD2RmjKAubdEvcblhwns
EBFqMLJfwOc6o20AQRRtYB8GTGTXBEie3GpY50n+9moiNMdimmBKQKBQJcmK2VdgOdN1ECs8Wno3
4Aky3kiDSwTb85SRDu6fnLvgim4WJs6cJDl6X+TQSmX/jcFWwF7JgyOQ0jU9V8XiH4ED8M3njf0K
x9hSUmO50wY/hYJda+/Zz5Lt/F6Aq3aUf9O/vVfGbI5T7wFAoiyjA85I0Qs8ceIHxCAZCU+Dggw8
0AIDO6poQLWbDKm5rBchP1YsH408eVrZ4XXcXHkGENnuPHU4p4H+Mjrb1dBWLkrQuCym1a64JfqH
8s6B22JWbrxmd0gtW1BUV8a58Q69F8KpizjuHvoDDTNVgFZ1xX1Eb+CatQ1EiuAjOLDPm2D+SSy+
jtr9HilCqYMKEhZK6qQ2wY9SDg9mElag3CIz+eJ7/6f/N7Q2ZHF5R+EOmdRPm1za+xf1JcafpC2N
2C3DkV/Hjb3LjQKbkLsNuTuJTauYOWEzSNyeyqVbc5VkZs7leAIjIfN6mpQK1JcFcG44sY+6O2su
5ARxPc8voLMOrqWDNLBpdGXfmSr4+jvsgk7KWxwiiv+kGQEwb0IAZ0s/4R5btWI8LHx5z1Dw1Xx2
Jj2VY1yRK19OM+i5VFhA6oaSSJY6FZRUAc3xvEUUQAx7FjTjAd8WZm6rCQLx1jHP5sxVAji1P3XU
rd9m4LLcreF/opJjMjWeQ+dui0lAva6AGSIT/U8UtgL4jhYPo+cvm2CMggVWJzuoNmShcVPirSvE
Wti1ou3S0S24RU+afTOQXCXeP7Wu2/36W3UEw67Udp2XYZMsXVVDFzjd/+96H6MrnYePeJqHU9EG
NPDh9G5kfoWAVRNSJQDd01n4HrqIM/n31YBmw1VX+Z9VLQmGBRKhCqVSOIIU+rnmy+aOZza5Eefy
OUv5obu3+TQBsKNs2yxeJuWuW2j7KMX36CLTZh2Ct2MdZlshDrq7LAddC4vxQ+YZo3yS5nj3cfVn
YHLm2zDbTMeKj1EhyRdH1MWZxsN3S01WdO1/GlcUKNANApT5SwmupIv6d31DyZYofzA0APCF3xgb
8BFdBZCzFKFZO2mM7oFWT+17IacvFtTg6dt0BmcVZs+zmVyj+DvWrwf+Qw4qOEW6w6BH5vcOrfdi
v7shYUe9lYJusQKE/lkip/XMJsL0pttGBQo4rb+GGwTak2zCzQtjzAITJvtjhhPrem2vnrSMSuaP
+P5Sqc5uk3Ij3sZftPdDvnZd0R99N4/tx+qSBADnAzhownZP+zbfnE6zcuHM/D9pz+OY3eOGWUbU
SpHqFNsGQLvOUQ6dBqWDeeLyylNuzInMY54XBMeDu9C9cJIdcGjVTBxZzn4VCBQxdWXHIe75CEWS
0gXnrAiRSZwON2099JPueFSZvNKwntxD8PV/SOvHgZBFrKUafsHN7QBjBWMMZHNdiG6wIjc4hmSY
P8g+8P6bRUi/ktsdiq1D6a56uK8KjOc4YkK+aX+TL/t7dxGTG3PP1+ShZ7mzCL3XL4MLSorwJcr3
rMpvX5Vd3l/QDGkms0Ex/MxbxFHQWuQ3Y7VzBhqrOWICUDTgBVxHRTLM1Gt7gH303rcbV4gvvxWM
7oyEVowhJHPeA3zQyafgrPzJRIpwplixBIcRu/vVNP4/KdhIJ6NbiG/uxZaJYlJ6eRlOS/np+BgV
TblHbEa6XuSAVmP1t64b8W004uukj9+z2OTfiytyX+ytdhoigTKuXXNmhh0gMlue6nfEYIMxyEhP
hUs05nS7v2Hb6FQ6RJYyX+IA0QcsDtfk8dJwPKcf2wPUtLa5zzjm3vtrKLj534YCmIi2gEQGgGgG
olY5FeH6uCcyqFz0EybORY7Iq3KeXelt0nkoHhmB6kXRQ5gaiqb7umSyFnfb1i3KGPTrUNjb04em
EETUSRWKwLEqR3YAO005cVDCzmH+tvPLQ8UH0EtcHYA1y0Uklz3W4vo19ko9yeUMxVG0UksgM88q
9RAG1iNYvP8fcifFfcFGiiv7VuMSQNhWxFQYA2Wr5jJsjkhZhkRj8oLnC1xkN0xj/2Oyjr2ieeP+
9uvz6oGVRxhz25SqNG1qjSkLJTKw9x6w8GwtVIgsR18u3PENHZsjVS0jHxlRnPQCyxNBhrb80rEp
7pkqoYoAvcG4jqnyc27pIeqykQOJdThZupVi+13ggWqzVvZF8pgZfLclUBZFnitoAZRQZNdDj20l
+kiXpaIGhgNrNLlyVCFWhZVmnIp8J7rqxiXo1FdTSkDd+aaTibTk3WaKfwmb+skiFHKh5zf254Ev
Q5q6Z6VBOHQOcYoPoRD5KOUT1fBqvkAXpuOEoMb6DBT36l/TW2RFp86Vjn6JVe5HqRJlU59Si3jB
0TnFgb2lLYSVKF9X5+uH65VikW/TzvB6vT11IxHrSa9YFgJMmKy/nbi1uC4K0eS8fTfPqbjUWBM5
Lw4fL/eGO0xsBaIYfPLsDyert4BUQlGCwKekUNgNNV2YhS3jnXabGv0VWLkZ+iVTnO3307lYY/ED
fQ3DPdU+82fnpJ1aSPjxKaPm6pEgoIMBQ7YntBDig12B2sSaY3Onj6wBXIkhOSbFvMjzbw5mqksr
roG8eoO6QKDOrcJxRktwR14UCvJUnPZxTeUR89uHQrL+TzFWfibncnL6rk3vrIh9YR+6OyOPph8p
s6224+uaImrJ5Ebju7jcHTQELREYFZ7NTOU+tSzQno9wNEEXlJPOw/T3M4NPb2gftd3JMt3ogqum
lGyy9oSte2yHnFO7jhGkt/mLogvF2Mi1JWjqmx9TgNVhnGkFgdWJP+PZ+WKqsBmx/fDz4yujcfbs
eh15vOr5fCJrwed9iUMo2yeBB6qZug43pCPwSUyR/f1rYWST5hsB/rIu0/hqOgJGk5I3ExIkr9QY
p2LFPY3moI2r1pj4V26Q8vigP7teU7CSC+Dro65PWHLbLbBeo3NILl8P3q7fX3TFmHjggUrQ9BYB
0A5k/R4ABwxw3ggZK1jEDQuTIrM25k1cfKS+asAY4280b11wYRRrsv+wlZXqGW/twFqqFBqxMdeI
ohyFTc/dfVFcol69niZAt1Lbpyouc2fUol9UeqaQ2xHDIePYLjJNSQ5cIiyIAYDL5L8QeVNOE5SK
4AeehhBm1s7KEX5ffJzssYu9GMR03f17qpGeZE2/wuAwytIHsb/yswifKaXVEwwb7YZaw8ckhbpG
Sj+S7SAguiK7OR34R48QXVIPRTSJdWB21ffr4c2SS0S9/+Nz6Q6m4fH4+9+uLUdVkO2qJvdVQFVk
LylLuKae+BRRozdDAnsTUhPy3PWat0rGu7pfG00BZ8EjyA/hrNJjCkAd7YmnMV+3wMTkXZFVJqxJ
kLS8fNZzbpVcDuB11OHgfxailr14ypHX0mrT5Wqa1etL3+IV/D2lV6S9tdDixJ3FlMuEdyvnw1v0
Xrm/+WpI/KMrsK8+mgl70pUmBo1QZ2jtcu/pF4UqpYkHkr+JPhP92aS4DM4ZvcbvhlKbOwE3UUDe
lKgfbyH3atnnWQ/Jvw6jfcIkN/P+Jm3VCI902VY/bG9d9IR/DD0hJIsB9WzY2qHzzjmfBiph0yru
A5nfh01YMhHTeEtex9AJGb3ytlBfqkSj7F5WinVgq8II+hrvF/lf+2qMS8GmF8pbgrZI1XWmsuJv
JeYSH5wHMWGx7GAzBSAT/lMHvJtmg8ZeoJ+Ek3i9pzddso235GY3Nb6AYSVIeiH+rZaRYFCWUk4F
XXBPeDS6ZavbTTKDifuBY/W9hvgRMwQrv9gSc4SBRVRU+cgHKrCOI7X4IYuc7hShElXWXsxhsiuC
S3b83MveeRPiDwTAIDgju6N9neSuAuyv7DIL0ZHnLfm9gHnqvZ9AC8MTenqMn4FPuR28T3nLnuas
+4j+Zms1VR7AABo3nTe9flPTvsq2TT+LdD/fqmpMHpHfjR8uf/g0nXa41XB2xgIbDmErbgfVz3WW
LVywzJrCm8lQtuE+3yv5CmmaTMjyuLMHruSAsMDjFKkcFbqzcTRtsexkjGdSFoBavl5l/S2SDizb
kY8ZZkKl6YIsAg4qFUvJOdU3RazJ7KmyjD0gNWUF/XoVJ9OIYbLXycHzUjsaKnx4bZe3sLUmJ5UR
3e1WlC77hdTC5J6TF7sG6ORdShA+yQYMkydk9FpxwCOHKrb7XIEd3rzw7E1+mRLUi9udvYlAjchQ
Mbk7cUDDBvn8/ZwOxJKcGWfQlXk07RZpYZV9i1PyXGsWxvQCgM4xpthY14PdpvWdvAfqsGpPDWHU
5PQ+zfcivRwygSv9KsD2vNTpaW56TuVLvTYNfzqIFidBfM9AC3HfhO/+d/TrF4zyuf9UPDGmbICt
2IwdIB56OPNBRwMMdaIsur7+hfx0kh/eVljlqW14b9V22gOuQNQLnwbn9/uBoiSh1TfSA0rTcjCD
d1dNzQtvZVL7cx50OUMQ/wWJH+JY9H68ztfS+j0tfDGhKTGytTt+RfpLbuEjRqfC4G13aEzZVFIO
panSszHU2WEwQwDr0svNwBVXp13K3yEB73bucsCGaHj5VHjQ66zG1Yl/jxmXsW27UKJ9wGw4unZc
/449EJtSSXk+JdzGbzhHYJ2hDuugT3sMNallp71nmU/xHkB6n6HY611swwlQjhYOoia1gD+uhMeQ
rNEclRgMgQcxqvPw0na1jNimUcv39clZuedgglswScBHbdfxz4U+rvR9Wpe/5wPLA2QYOHNjH198
DT+krv6J3/09oZIwdZYszaL51EOdw7YP2rFAyl/rK4wjCRweI6TnRo2DZu55fHiSYCd3XCwR9pi0
FtM+B7+14d2cwvfQEgVkiR3N03t8VEbUwmIQWBUJ19/6Fe7/VvfOtX7huc1aINwE7HNQ9YgIulBb
Hat8e3RqCb6bqNZ6HT/i5RdlD3psIfbl0uvkag0CtYTHLFMJD6HydKqBCEQP1wxc9ZwoN8FVtQlR
iPWjVKW/RFJH05bBgh4iFYOApO4eveYFOxymdtBxyPNhDHW/v9JSmHfC6CG/xtBWXpFBFpo7IW29
v9FxDKcFUuXb0P58VIC9tNfzNb69zSh4gXkSbRtn2QxhvODvHgwRWBwcvHSx00z0pa475DmDltoz
JF7A//rGI2D+5BWxvyFEVj6aJyufK2WmcWRFdaUn+hpDTvsUavgtDxNgQ8w2sTIPu1C+Vl7XUAGf
GDG2qkf+/CdTYWaRnZB8gwuAxPO+FgA+MJBaCqXJSeKEGQgC3fKIpP6UWTug0YOzmSsgFTvwMbK+
/3+9KliKRQ8gMXMU8tip0Dl8hfA8lImJidD1E0K4AFtXAxAZsoKPHKfcBBmLrXHuwgonazKCu7d3
n1GI0kjVC6Pvwb0fd4A9B3VkKcxZZvEIAJelPq/Wq0k6BDq8uSY4E/QwQQvCb4d/shCawxc3Dsaf
BhPxiM3RMw0EyFKGJPupOSDO2SPd0o6CK4UKGXqwJzoFd8b1dkVaQLrFjpyRkb9kHtoiPE9OLR2J
r140JYH7ttmsmHjqELbCx2S8v1fvK1wMcPastB8D4RK5FmXupAZamGUhw2odiSe+RP8hrXWEU6FI
1IfMROY7sMxXfi8KNluS4ipStK1eOsGoMGkMmTab2YygIc0IogqXna/E/8MHdDByNwHqqXkodxUz
WTRsOSEQ0Wzfn0rYeTOuxvc8NyAEMwhcgfXZhuLn5ScMTheqXH7aCbHY6AjXP8F4syKSOVa1I9bl
3qkKmxk16p5XMhBSzVbumorPS88LutcguOg/kbj45wmpN67+l3byuKWdcxLnoVW3o8+UTVLCmZs7
CbaLCK4AY6o7OenVz42w6Ju9k028bWZpwjUr6JQgC/omvNgVLdPkKyuHQ27ewToOotxuumsY5Wxw
7igMR+2D6kkdxYg6TxQmZVq6Jb3kIs8sTra9ziCxwgQb9FtuT5KFHNuNy0+pr7/WrNMG6/PLMvGw
7qcb7dl8GaY0fU6I6lgz5nr63jHdWp5JlwqxYBrvkYlaLk3oAytuQ0nzzJHxULYX4JDSF27tbw8d
cea6sVoaRmcx3DW78MioknSZYzNGDLcRkb7B9q23YRsQD8ayPOU3+sFNp1CDqFvmnUsUXBHjwFnf
dyJ15dxgxWkpz0QSExoogocrNQq7YaO9a7hEjMvHZoK4y2ryE+D8wUBRuSrJ1sTT0SFO8sB0g/HM
3NooSPbViUEbU99kcqIgsL1TAwAFvNoiz1DwC/vs+Z3CQpWQxfRz1+x9jzuB1wld2ggqMjKeekf6
8DHblS5J6RI6BWmTJZQ4ucncCgXdxuSHsszEfzq/dFoP5etopzrPpfmsDGPphkBCrcBFb+kEmJZN
mF/KJrKDGlDOZEP4uv05wLFVLF6RIUlufZkUHWJ0Kw/VUtKHqBUKiuUR7vq8O2qLVy3oWZbwZKUY
82i+fplIoe3Ld8mpBRYNtx6T2eRsLVRxhVbtem1fqRR8vLuiI7D5yJU6oI0vYm7HQTbFj9wd/5dh
H+S2Az/1JWpXVGWLFPLRbcCHPEG5cD2GDrfMn4Am457IV/qIR+lxTwB1VCZBcc1cXcedkM4sj64/
hw2Q4mRswUJlPc1rcCSssUHyyOXnlQ850NpZbS85uoboejz3WO+NzLF4d59Q1rzBPphaBVAXpH1D
KoU9uQ1GCcYmzxopJ4JDEX4uCu8e5uqDsALNZ9ppKlXNO0wMBiB2/rFSgbkhNbmcPrkoUAHsPHEz
BfzkawFL9OherI13wqzGLR3ckuRb007q4lkeKmJtUABuj7G1GWXsdD7AYWraHMnOQBdfdrUxL8Vx
Qw6+S7HJyR/JAKtK0NFAaogHxz43FwSWk0LPN4+7r6G0SF9BfPImAsKh+pu8eem3zl0/4Kf2OFIR
tVA6hbZrGDmrULECdYyLQhLZnH9TxEdElO45La4VFK+7Skc5va0ybwkWfnWLrFDKkYR3SDdgefna
HCOHCZe2AalZDphLHcrgZ5nBkyrtv2koXzGZ0Lw6uQbf5bv/psxdVvwNa91c1EZ2yD/30u3DSYtm
SnEU+lbDrtMUIZRILzIIsBujY2M2rwm4QG1mS+CY63xQkvL8OvBffyCqepdRh7hp3SUHSsDCxLKM
klCWeJqW1/Ba1+0zhoAT7rxtfmqePRbUmxnv7se+Au8ZYWUW/F9iFM4PqZiMoUbcZ6bdVO+crdL+
RxZ15RmLahBlSTocFuTnj6mC2c5RmwRInt3Awoqr9t292x2C9V7oLJpsILW63yr5C8pvlVLGfVWV
dHXW2pf5JIwp/zJ+jx2MzY9kALmBuHdGGw/BlfAykOMt6NQdKrIDyK0qOLhIg9aKmKkHNpbNdnS3
VOnbvVOmmYFxMjXJtbjEZ1mRL7HbXiiAMykBam3ahnlHCft614TUIyEdIDd0MopdO62DhTT14WRx
1Oa7V7c6rvxJ0BBaQEqZ2aVXgc7ubrCBCeBIfUTVuv99Ev5qMvoyEOrzF60IjmTN82MKDHIamHZy
NM7AvUcg8UP8j86IH0znaswYkmO2tszL2+10t0iz6GuopOPLu4iau6w9Kv9/sZAY1x+yxrAci7b7
45dkF2At7vWaUF2dsk7Sk8B8Jop1BYzR7jopOCPPOcQLzmRTIrdBNY32Lxl++lBaTJZQf9/MhDb3
UVOWb33WjV8GpMq+aSaWR9oIYcGjBh9LCbN8mCfsAFGxcadi8K3CAWh69BgXNnoy9nAtGu2OuTcO
RkhEVvaGaAsgvl4Rrb3jKjXRBApQZ4tNufSwMDP6dgCo/GGcGoVG30yurhgVmRlwJXhc9w2XAt6T
SPZ7Bx2PmfF6IVweW/2qI87wHGp2PyywBK2OTK91sCqCwU+jQqzgeGDmSBnPtof2QG/0bC29CdLt
WL6H7Z16jDUATAvVKit7K3yXTOqWOxPHbl5+Nf9JRRK6vZ77G7ITbWWhb3Nv3btNqI45N0Gp916j
e42OO3oagzznznXtQUwYVfKepgiJ0N/uttEuLlFpagsKcrrKixSPbpsA1lGBmu1fPdzFSYdG4IIg
guXuKpzisToILphCKCAsS1nEi6DPOeXOdX+NKRMaciLPXlKHUA0gDlnqGx8WcNJKFX4TMwv78pUC
aFZi1bIv2kGVX67nqrN+7hiKr+vSl/KPbLKXR+PJVHIMA6ZRoj3TOjOCC3p6yrSeFfGn+Y7iZX3+
zYqK/fSeBp2bKarhZygebtJ1fxBEeD7ULFWtaSvxX4baGeg2dwJZT8SWOzQuMaVcdekG+vVq3K81
To2soKqlchIqXNra8CLiheTjFRg3pIffjNokfvT1AtT+ZkB8w9jYlj/s7+jTzi12mwJWxl4qfQA4
Yb7eUK+nANuNSIH+91xsQXs/x+SLfGtlM2RXUH8mohN2X+FZNBCZ6EG6ZmyqSHC19+ZtW8AlzabE
1PG5d944/rKPqrO95kHV0/G6wamr2dICk37RXG/j20CGQ1bIpj6UAmSckwdtVmYBh8SG54VKkkQz
iWCJHQAwNWgv538dSS8Zi2s29BGOV946HY2p6DGKegXKwTG9eK56h2UxNYLXU0ZJhQUpmgt4g24n
YvgmCRGjh5COcUf7WY7X3X9719AmLYf/de74GX8QDELvphabevE/Qy3+5ZFpQs+5/RRpFqHOH8D0
z7U0mI4wptBFFSMZ3Ng80mKbolRABFj8Zco9cKN+m7/Mua07dq5wmuv+QXS/jORvrZnhDymmfTYX
jqD3PQ4aVoN4hSNujnYIyivkykAPsQPZT+8/pO/dxse1CacjLkwGFx5+Hedu79x5d6rCbaGpUfjF
Pdag0j7HOnRsXvNNPNiIb5TEXGP+VPnjl8szoOxWyxJE+jZmOqvrf5/RmrDSIUHX5dIXCP6Rh5qD
APWB7Y3SYZ55iITL56NF/Pxwk1rAzMAtw6x4E1vg5y3LYl4WMfU/4v9UhWXQ6AyPmd9I/5w5aQGO
AdinqYFRLZxPjQ09EAtP8baopIm0fE77cMw7fPa7iH22wPehK9QCC+1NuZxslNF9KZkQ4sFUCqu0
m9oe8LMEgAN9z7DDNSTpOO90eqhg6LbKsHgG12LnnwnjlhUI5Jw3g/OU1C/RJYjCGErm9uuaLV4A
IcMztgL4AZsBgXiI2wIaPYr24RkCCyI42kNln6nc41UXxVh4V4j07jSDc/COfVdF6KAla5w+CMVc
uzKXCXGn/ndS2GReAbUR84aCpcEZUdVuXEodBdCD4kn18sYefgW7TEYgRu1AHZ/uauPIhdrGfZL6
3IGL3wacw6rck1K6e/ypbXDisp6bQadfPyOqSmv9+d8M1OUw7obAB5uxmTkUF/tFDLLAX4iYMFiT
avscGQC/BzMuaLUkR3jNJHVFeZedD1+czLKht9ZKXveQrVbVEgVAca6CAJWBfkZMnMyAwf0pSVHl
VyVnz550f/cPEzv+dGMT53GmFc5H+FAns018bJXbJTqXAkpAWNU6fyDtHYDkiA7TOio1DLH2Dlfe
2UtfN78zInv+6YLdLTTnvYBT7yeWQHurjxMZZrogcrgX2c8j3tqmGuV1Op9zCeEG+S33MaC7lY4S
4fUK67oiHUjyq6FKZoNpi2FHN8dItyyPTWntINXehKrSPpT+Oyt6MA/eMgK8eQNp795Jry64U2Aq
qjhKe5Y5slfY5oV91FNLy1fFmtezqmxTPzWNuJIC8UUl8hsQsz3GeabgkFwlWAQClQ/kqwgjDhr1
Hn6+HCRaKqBSRWo2Z6I3Blo4lHG1QupLeqPmO50XW+/RbAkdAddtJPD6G1AjV9jXtzmtBOoo4eJe
Tw+R8ajfpM54LSqMraX25d9WPmsc98mPXG5cQ7qdJ1tozX+Q13yRtEkLMw0YDbKbgbOjR9vrlX4B
ENSUF3OYxgzKx4mTuFkdi/bi5MsqXYO8uYj3JLudJIY6R8X3DMjOBydb74+xb1vB/WoWxKwzZ1Ah
nDK6SJymunhUWFBB8Pg23dn4BNm69DJwX4f28z0W9QnW4QzEuqG+Swl/GJxcfLluAnPNPvCZ8xC4
cWuVq/+FYJKAgB5hGv7M9YdMTtzfI08uKdB+BV+AeogwYMElMvQU9eSCdg3A3pfgOzm18N7CZgUu
JRkXH0okgYRa3RZnXR2JAFlYVq0yEl45G3Fki8dkGtMMP4ab1gIZwK5XVROcOMltLe5DD2nhsUR8
N4LNs/fLyNuX3SZjxNNTQA06wFWhL0qjd4phQYHNLa50JvoSpXNByeYgkmep+qDHfrG54Kzc3wou
e7ITe1QaD+gWpUzC5doXhChonUvnM8yq+BXV3KuHio9HL9wt7vlMci+VaDCrWs05xvAyTUMUGGIq
VNRW9BLUv9bj8vkcBL2V4Xf0CiNNGrgsNzbC1bbw26yZqlcto58+cVzhMqt5TYJUq1Pjn/GAQauZ
7Kho4n+FKINXUSKLwg1ZcACXEO5t0afsi5eKHGB1D/k17Bjy5yAtFD6VJhNhjtBg71umGi3ZLCwu
nu10F4/uZrSa0NufZiRJqE0Ya7usXqdkF/EFWl6n9wUSf5bzDn0nCwJGKjqMH3PjKvPuZul4Nm8Y
wYYTzUggG7uIG2OzA/+fdorsrmdD7YqBScpOBj/UmEMPlNZPUPZodSFZfFE0iUGEa2Y5w8VYwH3j
JwnWRxEwn1mUBUOEAtGE+HUFrnHncy+R5ehxIjP1iqYSmRuK8XB1XnUjXy6Un8H6+YlvyVNV5Tuf
ljf8zGkEYIUXBXtw/VDh5B1NhyobwAtCz4g6cINfIKTPyH+5+p+fzyI/6MDqu7Uj6V3iI9HrBIb3
KWnGNNvlvKKF112Vhdo7AYBVAF6AQemtHmePkpOD5ar4eIBYV2OIsigxiU1dcLvyS3+I8OGFwJXl
OGTKXeeSVCInywmDrBlBJpc/B68zOdkZ6MWo3BVyT0Eceja38zrzFuqFBuL5eleMFnWdt+zc+VnP
103LxdYDH2/RY7byuQhAdbpzlaYntKEUOh2vAW6b4N5yAo4GLoAM+LrL+uYA2ThYCD93evRRDLDj
CCYmfKN3nvbjnvMqP3CHAHQ9F8kAdIBii+OCgPtb0WpZlAwbPDaeRolp/oenuIcUXTYyLVX5JrFB
uDnL2W8iMjJNC+6Vikchmowbfuqfcqfto6AYhGaW/UyPXC/EIkOQEuMwAvRZoldvLN1U5MG6DBkp
41po46rz9cE8LdFbe+gz8u2bKyOttrIT2/D4bNqoqux0zfY40re3Ik62cWpJhosEHKBJPP4Yrxty
h/D2SqRYVA3TuJED+qgo81E/qWQRtwwveJCsNgrTDta12+fIMgO50Zy6iQMLKS8olNMAA6LplvmU
pERAVqqHJmPEose5unKBldacHx2HxEgnCdJ3u3cVVPN+k9Hhfg6pq5ZzpogDXodymZMPMwV1/Gi4
FcTXEo9ZNoBQwjKBRqSkTPlzh7T31e1ATsTKU2TQYf+z2fTg4+cWni9ZuklQQ8y361Dd8g/9gQmm
rAjyEStjagnYP0dQ50avkFyDDy0GAKQfPNSh7n1OabjGPpT0J7X/Vq1ixDULCO6YWqJNpYuGRM6R
dJAjNfiAmU5HjP0Xf/q+8c9+l4Fo2xj6vMKbNBILD+oZ38IBWDOs3QFbZ4ir/L8XAarUtTHuKrrH
Qmxe1WXnz5vIxFc5H8fwEgRP0UWjeJbRK6UJrJ20B/nlaITMofrNInpA58EebPvT5rKiuQd4KCNg
x0diUCcYl9UaUqzOTBCps0wwei+iwsO7DMzhC7GN8jKzkqm41w1dCHXdLB0EynIk8TWHmy1Cxr2h
c/WefpcJzh0rBNWPdICiq1hSrJDEjK89ZSlUz69kQYuhNSNRr0+JZAlrneqvAq346KjJ7L31gAQw
WJ0+Rf29Tn/rbQBM3X/xHconMfMi/9UpaqmlxJXw9kwAuTrUw9dT0NFRCqOU0OPZAVhmYm+NIMfW
CpkJehQJ4AIm9FwlXCvsCWpaYRZWGaBm5EfE4xm4K5flQP6EVJp8XJ/jyuXSV/Gt+UUeGw1852pz
ETbhX/98ZSEvVEVzAl99tHZ9ecBYhafyOOPc+I7/tra7UlbXt9n1dOu/9QNdv9czREDtoDLJPfzf
q1pDwjpK38+qWubAjwKJteBX242bgh/URSGWD4UnDdNEZpp3E1CMce7BofumEYv0h8a3/5ZEF2uL
FYwL492y7lcxq7O2WiBFgQYKIHr0X244dm/0aa3rLnKwMk4UcVQZ+ulCMi1DK1/CpP4jByR/ZSuz
UCp19zgXxra3nzfzO4T0ZB2TMMDOVoAk/l6j5Zo3q/FKgPde4D8hk3IdQBmpQ/PBj+6VviOofY1j
Uhxmg/Od+e2IT2pWXCvO5q4ixnu9g9Wgqh33WrmTyGxEKf0NS7/Qt5JtLEngqjsoJD1C3wTf/LM4
99qyFyN0IP7kfaUbco7HPEimsprHK2rYqcjriZ2x4nNo88l0/VDaJwWo+ShcBnpYMuc3H4xutxVf
gJM+UVQNuiXrAM/MV/jXbBMUPrZCbDVLIH0jHdnXxmIMvQ8g3xJugAqs3g3Y/4m6BKHRz1XHsYX+
ARuOJ0LpK3FWGRGmz09xVLiPFqWIMCYztm+9Q6w8shEoTPbsx1e6O8wv0Kmb7kQKTHCx5j8IehcJ
U5q378wa5e6/Oa9M1iTEM97AGvnM6C4CSklz36VNshJqQ5XQRzWB6zaEeh5bQjO+NZ+lXaT2iXRJ
IVjNpmgxkr+cnt+bNj89HFH1+sSExrs6pZyakDwqwDA8ZRqDce7t3/qt3DFup6ohceW+THJO7GMI
uKJ4D6gcifrEeH9WB8Z2Ye/D97c1gwadky8aTvATssUElHWs9td5nuI01HbcblauS3o+xDBxvoX9
n4nwD/FIqMi+7yifOuxVf3HHoL18qvmn0pZhZL9CqMxu8P7ls42Ap4jvoFw0lZMSN8m5cuXG6LDR
Scn02iuvHu26AUyJ+uIti3x7YcEVwGpzy3WGoxkDq8ao/co208kvFMJn3fYhI7q2W5iI6mXxcHER
RFspOFQJCiAmTWB6/nC5JNCiV8YQf6xag0jYue46VWnkscUx6MLM/aOQ0+w0EXLLQlkgba6MGm7M
agc2CSwiMpkhKOugBy+3aGaS+QdL5tDkreztn/WyXvQnF23pD4GfeRlZhsnp3Zu/iGGDDDk2SYpB
N2YwjhZhkLTWWLShl2hYu3bCjcqVAIFfrPobPBqjHfyh3y+Eu4xfmT2mXM67EwFY3Rm2ATtC/7qo
J3aZ27kx1SU0YcgkwR3d3mDqX3Ww7dZp6PTBjn9GQsD6jDwrbxBkk2sSDdtko54miaPn6EwvkJdU
AYgFKMY//nrN9RMKCzehSrIQXy6czv3wp/9IfTcXDcRT1K6h4jnMkoQ8NXN1RaR4vJsjWVjyfG8x
+VXMUqXm4Y2tf2p27Nm3UNzLYW4ikFvh5Y2+ea1IIkIszMGikIHVMm9aR4wMcbHZNZOw7zdhZvs9
eOUfQR1kZ9uDm8kqmw15imTW5B4gVRXlrOCsvw46JWi/ioDpRAn3sEANiX81/NUS+6RSkgLyj8sT
upQmhcYJvW2jpKuvc5jbGLao72c15bYxIsSib+l9DJJf0Y6LJ5lG3Iepsp4Kn1H4r3srDnMHrZYJ
VHBzT7P8b43IwKOaopTvCWkRfkWN2e+FkORGKl7RA4Y6F3beQAqoWCIBHzRz+lMs2PsJllOPNDJs
wI+a1QOG8MdnmwfUhInj9DayZiql4KZUJcy8UChbVteaCT8FYYmDaUGD5uzbnnVEIMA7BJPrYc7n
yPn8+60hN2NcoYsah/G8mvDu42R/aqgGRVArN63yi/LNBXFB3tV2mmk9KWqeJpUPr+kljdM3Y6PV
uaMzTMyY4dUAsesh2xtMC0gXMUvmPL63ibZ1zJDcNEN8bivu18aRyrSvxzKWpta2auXFiFOQNg5y
1wFxDggGqc0HVuFG6kEjEON6YTO0l+4/PEnTj8G6sT/Ugfd0HJ5HszMT1Q70Sum7SZCO3ZUrMH8q
Fa2rhIiszzzGC+BGSNla4TE8EFsnZDttMJCY9rn11Gn7fETIsb1LQRoshTJ2U3+/vK+caYe1dzuU
RaBdTWjUoC6UYIGdqGmAABgLmQtUTQ83l2vkQL7v0F3HUC6ym92peKZ96tTAruzMDj/d+pIXrGos
NfTEN0XlKZfAHRXdpzPKQ2XnsOQeB6HJ9MSeKpTlVXcgHchgewTF/MogQqck9hwSDwMAa1ZXzY8j
iwKhEu0ZYUyTSK5s2oc/ajWcFJfmlBwlADVxW56AsoEUn0tLTxx+knYOh/7gg+24ElXQn40rb3fI
l+Eu0+/18XzQwEDydKjNSQIUBo4PBfl/apIPWGuWVE0uzi1Iu+zu3dtveH8ZzOwOOzwY1zIm2TPC
0eNFxUnzR3iJ7rR1euOzLyTXCHiygmO/ZPUdE7e2kOTvHY7YpxJfPcidoLQHDey4ie6nt8qMWOdw
LR78k/qJnzNNHohNJTq/h0s8wyoBDyLMZITsXvFv28Tx9GuUEjO++titygX3lan3nkxNWmnOIJVe
+iC17oLdMOr+/kixupAwUvZPlA9HmQdFMdOubWFcXB7ICeHYtUnZShMoX6wMihEKZRHkFB0dFiE3
sYPYO9+Uw2tScnYxQX4UnBZdry/HjziCKd3E8nh+5NG8tmfOXsP7VOtsqh6qIX5uei3207yoN56+
rRE4oaTl9ZZzsIBooyYh0UiVVyqTpvB+QlsFnJ86q5vCyxf6BsEupyM+Iyxhx17+6F62MarwZLZ2
UlGTh4LCpDJML+63el0YRHGVWEYQBt2ZS7DUa8I/X6K5FM4MIIJC0lYAGfXKkTnVYqewyf3AZy7Z
HHfitX7w1N2YE0GGiCZZiJtBrBS4U++OcnFwSyzZYvYoCj00ZPmfXqSxAfMd1QwR2E3kUSWL2C9t
3aERPuMAVEW1qcrvENkgGBNUADSjc2PIgV0hG/zNgGf1HVFsvkULiaOs8LrnkusXU0TU2euIXNIT
6MxPP3TSRPrWT441e2REaz1S4zqBmnvqyyXUMg/oqmhaJNXAjw+cAWFwK7H1v25D5IxfTaRFypu+
0uFDUW5EMmKHvdUZDaifG01vyo7XJFO0bVwkz/1XnBLqYSkgW379odVMrM/5JFNrwHspXF4CN/NE
Bc87n2wk0hFmu5+hDXd8xxvMitVv4ziG+0SfUwL9Qr32q3xjVaJICeRtutHkcZHF97htGD56YE0v
gJ902AhJp8mwpeHJEz0Zvu5e6UD2QvaD5FXZaf/fsxcuWJoJwcmbYJe/lphwIeb9tzEG9XolpLuA
R8S09zb3yFtINe36Vou+Glpy/mcbKqQFpqxqsC++C4+JGEPkU1YnoW/nZs2wzcn0/kboV3fukm+h
7sV/hg+AmGKbeVCmQ9Le/mQ4NVQSYb4605cN4KkswTD3660A2+yw3777WTbdfRArRz2ERqA/bpEZ
Er4PtE1Wl2nTOXRPOVqT55JmbHuo/zMnxDDIp/MqyHTLF3tRKr7Mqqo5HomuX+MMeKhVfjmHDX4i
3Cgm9XuYdTOxLLdOJxJpHUTT1FGmQef60cjphnp0rLlAamKkqf9q3qOCbbyqKu6CBnOiglPvMN5C
Y45V+OAxeHrbr/CIIDu4LitBQYANUISqlxPcFt4rH0WHDy9IV+7cpH4wk5r/LIQjHa0kkiE3hvQo
hPM+pme7Y8v+TmkFaextLFG31Dl9a3jDOlmNOo4vURmsVBmOJvlKcwlg8xTBYCj4tU/4qAsN/FEE
eO/Mjx3TmC4/pH4xnucYgttMcRnpYzoHGY/VwZU/0SdGBQKmcyvDl+Fz43MKPAhm4nP/1ClxU6oJ
7TE7fp0LTpFzncnWYQpZFBX+NibrcUP2tnxiCUjyTemcTUxUUgMaDw2RMBLjGI37rRoUyX96kAX/
+eRuwdvVPJrY0uB94ZdFi0NukqtJDOTWM7FsbMqrK9yehwUkuZq3cd7mvSG6imKjBkTwqRST+6Rr
qH7OgytNnB9bERRTeLByVPnsIg0FGkBkzxYNwTyZFa6quFwRZ9pjFzJ32mwcKlP8aNUFoA4ebhaY
mjDx33OI7gBMrlA950mcvH7i+rGx5QZF6blBLfXruBLebK6Q4sGz1oJvIec3bY41VtAOwH7hOYem
VqLMWQT/OYd51twFqScDSm1imKvLdqvOOF8swqZnDk06FL4S9I0MBg3VxgRuj+Cmupz7uUDLvDdb
LF+a7bDYPIgZv6fCKVbbFww10mDyFQsKydYkdr/7/DaJk3bSr6bbfC5U4FCtI4AcqkxaVMIvEs03
eg2sT46R9zJ1fb4AkR+k4m8WZ1Om+QzubzwPGHOcwh+qMGjRpDX/PVMBnddOjtnOYFQiSVWnNvKi
635NCVLu6f/Gq0cS5CclK869Pto9SlxMy3sMnWhFjPySh3ljugvGT6zsOBjGK0ALB76t6r7kZq23
bWS4GZEFOHgAB6Il1T1KBSQx1kCvRCs3CNgcUBd09PH64MDAuyAysP+deExZGxLTevRONP2FTxIF
JjxPTkM8Qo1PWJydACMwTy1a6Ps1shtYNY5XQ41js0p8M+8TbGJYosS0uoOpKQrpObxAJ3M7NMvN
EfrEp0GW9QtlRRzbPipw2sO5xwftOtvhEYeJ4k/GQuKaOoc10UU1POtK5fkLgEdEjo1CHwd5hXVV
D2je2PjY075PDw+qNJTAYzAWJ9Yvhj0kkcYdrA3iNoJOWOUhrX5PnBMulUp3im6TBLWwCVDIQTiZ
7yzuvrSA6Gh3NyX7wua4YeoTRg95shlBXoVvFU4Tj7/8qIG/tG6FTDoqZLgxLe5RnFM/Uo76LZFI
4pkmp6M2bFf/F1FOIRemLgisPJwWz6tSsag1lQSiA7M8G19CxSH4EyyEXC7Z8yztnmGLFiwFnhPn
8OakVRl7znVxqYE2/+P004Txj8k3yBj+SU0/xCHdOeBmoxrYZ4U2Ws+3R4ZUyyPU8wAqepGR6dsE
SIIG1GZ7G60uVTt6o5d4oPJAMVdiWz/KWyGnifujlKTwjUWysJdNBsF5CEGwur8QVJbhzWaWYWtg
k69lPBrkhvI3guzuVmAzIxMqioJqUneo7d02PVTfrEm6tUEI8a8zT3+2nscNRiQzDnm4IJRkeeHF
oOpbZ5f/Rt/wv7Sdls78uvExGN5rC9tgMdlSs9nTFl7jBtZB6AIlxpg0AcMpiohnr0+k5OQM1sEc
xYqVQYcHuGmq76Ghj5uWuyIjT/4tIOuKKyZrHd50KVN3+yYumFzJi3tCY0owwcNz/RGRDUTHEGZA
CNU3OGBzDZ4kUQq4JQSMY3qL16BjXq6g+RT0lQs1jjyizYWN85oT/T5wwvZj+7zpchT0/uM1cTMl
9YPQKHI8B+5lPpYZ0UR43uqREUY50dGrECfrgyFYEmmLRWMF7Tj1FOZ+2kriqPGi/L3Kja0tOHPB
KwHQpKJWbS1zQReTjuCbQ/UB1eIajgYnUQPxSHVhSi4AfcPoDe6OyFmw9g1kdTMAvNIP2OV4RPYj
U6C/0JjVaJn+Iz4P/9meDGRQKtcr1EUt6OUGq1Cz9kbkXL1VpuI9lXASB0vyQfkUDhNk+zlvqkHO
BaMtNiomCNKFerkYGpiB1SagQKRiDwikX+EyeMsW2l7ZzNmlhjHy3BdW69TYTO84+5Gy5R7nzIq9
k39L6DlrfW4Oo6EQPHsLtv7dBmbSwTycNuDtT2js49sw4AMnCNwWrdAuEH8ius0k9lZ7EaEKkJBQ
EiaCx8RpiFe9NXPRSGE4OnXRMQ1ZjsbosBEIyzNDENtRyZVe1V1vECUGL5HpgT9ApNqHXpB8G2FU
Vppg/PiPEYhYlSSHcdm78iEaXIh2LT0mzDQF5ml5JNMCbfa4FKtm8zpmuSBwSkHxktbi0sVurgKv
NsgIHcbMDEKR/7yIDpP7ZyJsMFqs9NLUk5BlZjn/oZ3UJvCDP0xnDyaQU294Hfjbtz3FAogvLiRY
/QZ2WpvZKCkjJcEwzxBHT9JlGLd6gvNxj3k+cxLY1jLQZTH+yYJcpTwHbRXsFt6iFkQdOQuWEfoM
RIrkm7xAsc5Cu3GafDFdFjwlSgarG1cNPhOoENC+AmBuCPNpMdEUnoh/Ar9wzwjXc/ymGbOR+0RQ
qI3dCHvdF81B0WH3hx0+qLDoYG63gmWmNhyVVta+WvsVK2U3IR6cJt+Vhjh9HU3QY/D9HMTccaXi
SnBxjJMsMkKvZQ2XBQ3gRxIg7Y0gB5P+diAr1vgOKUGiWYb7Cf/MBkmTm5wEhQZ5a8MfnyPfcX3p
7jOH10vKmMAyZDNXzpqYF3Wq3rI+1cpZWMWe30TWBj5WWzzH0zHZZ/Gqc0tH0vzgAQYFv2qrQZdN
sge3BxdhPw3uIAeUGrw5Of6yAZUeVZ/y67XiGwhygYe7KHblzaELNtB+j957xZfrj4fkMwiYJGLA
wrAQnSDdQpxK5eS7c5nLv+WfjS0bdkEMRsLe/66ndSmSbvch8tUNojytYD+y4ARJxEVeuifmTllw
lqAX8HV8Ao5zGX1H1xQeuPclPFSyjsIJE28dj3yEjoNPEI2824wIm8gMDScTz6IWrMqclsYYzl/k
74TKS6Og3J3lwtTWWflepTRxnndsRmkWAOmrKHEZ+9WF418g3Hmo2qNpodMaUV+N3sxGqgqCFkJb
LMBipgy8+Nu0+EM3uVh9Lq3bF68L+kWBFoJ8hrs3fV79F68FJ54oQGHLYf/5TnuQMZMWXJjJvYvJ
vx8BT+b6SamN73NWm/0T99EojA6lfNl4Ktejm3BBgCfJEnyMLdpKxNpLYueddrqXE51MRWk8ictF
xQrooSTSA+vM8bcRECMsscn0KFtgUrg7I/SLLfutmUO4oJMD+3P059XX1Y/FW4Cqk+kezBK6eA2Z
eVxsvtBt2H/O1LtJsAvncz34Ivl/QvRNBuRCaNy5nuxhvo1uV/2P2nYnK8uwC1Vdd9iaX6j5/n7t
tPYpGBa9BDQnMvCyaOrefgGqCynE6nhR8sV12Di4aIfIZ2nLvGdwcaxHONDJm44Ogqvf4v4MB/qI
pCK2W3cwrH+Y9hpaZI4SR0fFmRHvpU8hC985D6Zztw6XHOZVFP+XOrwqnZvV7k8JJ+6tc3SGjHX6
ohrmFNSLIzctXWAGDdqkTgcLFnDhva5EPHRDS7h3RKR745DfPnup1SOOSYqR9+tvI6Asj2M3jlbH
U4thDyt5zxOBg/7FUQpY2sPihd9fuHORjPOUOGDphcjVCvOFk+RmOymsvHbBv8gqwWbq2d1vLnGY
hhhyOgXWxYVtj3V8aV0aSqYlYWd/Uo6lFXlGpOPSzR7xHqtb1dtpw56vK8rZoiznISyEnwc3eNoF
8DxFLZi/lg90likt3RcE1al3wABK3rcKMaSNSxirzg1GpX+ARKA1B3Z2QhQYS7teyu1iCq9jUfoU
PZg66Bt5J+WHkuPTebaSlYXa8nuXeb+YtixBf9ttwephnQy5FjxrB0rP0/RJiHgVxjRxX4ywuW3M
ekpXzsWCiKs4N/5g/wk3KXL7TPVqjsYJ6lyn8BW1ukPoE4KHUonrZeJZs9fFK6MJs1CJkOf2+mKO
mEGevLAMGQmxtIS4tLTpBS7kUkNQMWWUbhmWCt7W2VAdDLM48DSqqNXgUwVoKnOrVJF5ud1TiiKA
QBYRc+cQA3zMDg4A86WYp2lQe+bUNtZDdWVcmwZJbVC/OJmTIbI9K/cQZj7KacngGNP+SV1LVacH
ObnwYLwjoYqbIB/Sc9avWlbvJmkvSo2hvf0+Nf1Ttd16SiOXyzlZoOcpmjoiXBzWin99UkxOukAh
qfUhgL51UnmWUz21z1oR6Pl4MuM7dkGMf5+Yb/jWcXYAkFQlUe8VUIfiI2K5U0ErcUyfUtRYxjia
Xj+KFLyi51LaER+bTpmJrANEp1QQFZm8Aq9bVmEwHoJ5baxicfLKBAlfXuxpoJRb+mxmFlAV/3qe
yF+spMejZfLr2uAWkiRNv6PIstGNVuxev+lUN/hFuYFJ4wLgHqmBiFIBcz4oy4t/i6hTseNRzcpd
0ihuoc45cGUfp9TtMgfWbP7L1SLb1aXwzfwZ9Td9pMtrjecogZa8dJi5cPRCdoR+fO76CkPyNTZa
BrfmGZD4cc9LfgiFkOxx4qDzOW5l07bR0IZscSKpILOkdvwAd5/JqKQMRYCHGMDp8MhIAzDOB15O
QnbAivopnGjd6iYZZK1EZjxanGKA5OX9JBv4vyuzHi3/O1GJGoZj4ZP05WlARi9VXUlTgCGs87YE
TLwYaHHoL2JyTolRU1dR0G//h73YVKqu8oPOVzQlu9ANMs8YWTPKNpjCPEE9sIQS+T0jggBHieoj
KOTnxgQELj9VdRoqOXUGXegR3X/BoIpL98s4N7nGVCBGRlSZ5pUVeZPTY492vQrujFVWEh0WP1wK
CdNWr05ftvhZltcWRqCGWeUyQSkN/FKXOpfPOVvN4aTbJxEV/8CkvtHIl8yPVYgclm8LcpJe83HP
k74Q/gbAwhbZK5t1vT9FfvNwHtkDGQgJxkaKkysXed8yQQwVDJpVYRjMsb0OO9ATtu+j0hxsSftA
bxoj3O7cycGui2F6FzFaEN1ytYLHVXoULhZUKneZj+7gIHT/3/Gfl1uLYi0CcCkuRvJwTqaJjgdG
JefL19US1/9byxTTa+gKJv4+ilnpCxmmB0hDnc6eWwWjlvjS7J96/IPXDdeYPQBZr8RAs4Aii2xE
ISy0lg8PZ3yWfcA3l8RodFB5pQNmsbTWiSHwhTBAqRjDdwTCfKTLzZC6EGq8ZuxZto0kMmFBrH+z
wQuE2Dm+5mov0qAVZz9ft5Hk5ESSzqdW+0wQqguAfvI00QsglyKl6P/qCJuvRx7neH4bJoMS1g0e
Dz0x5kSHYx2GxTaCF36cPcnDizU0jLbCTVn8SS9t4NFekDI9gRYtxCgcUn74Oh7QFBEcxt3hB3ha
mZlp0+2dKfGnBHL/nhDE+5+HCUPNpnOhWaM1l/SEpdI4OGopQqCFCjwG1ZeZqZUKB2Wq1yto01lQ
jSn9zeovstKK2jZwcoyxmngtH7WEOgLN2hQ3Gq/Y9fGxlJydze+oZBOUadiloFW+1wmxBQdJzk/0
94Vhv5s/c0l8hSKOUccZy+LBke0BMFEU7fOD8vdptd2K/n9Ke9Lh8abaCHa1MC8nC9mk7JynJiIU
xhHi2tuSyPskuMh7ICLGtOiPtdAGtVdn9Zy6M69+7ShjyZLpsmkuEJQBeNOYFPoM/1FiM7DN6DL4
qVj/Gc3aQnj4HJJCwR0DXifBeSFlW2LCiBGnh49EtRYAKaFTgW4NHTJqABKeO9Pxy/2kcf1RzSf5
RFhHiGwXczETP+1aNfTkPdm7np2/igZralA46nhtHtHrtpVcdD+ED6e6i8aERUJGDJ3F/VJ1Drz1
sTphBuOd5oUl1yBdn+OkMjyL6AJTxiBsU9ORRCNd05VmiI2qyb8t7SBtz6pqmMFNAingACvq+Bdv
J6FcjRhOFFMysUzMe0Tg/CWyyCEgNlBNJIACp+XegAaDparse83bh3CfYT5uL5QOGN4I8clXI0oa
8URfOwnvZSed/NUQnaD3waOtUmvn97S59t77aQAsB/vr7TgLrNk5xvVIomzvDCIY7HZtVoxNquPm
Ksst0LONxtPTFf2PCn9qw4z+XabggmN4CL0ybhfq2l4rKW77J8ahgQyKlbTYRPvZMI0eWxMV5hIM
hHMCGdIHAqG3GdQJyeosUQoklSN+vaVRNuuGk1TNm5yhbonP1z3Njd/b5S9Sd0d/DU53TReNY07F
5iFiB8clz13LtCPb4/vh5+sUkuWONG2qDlAPBJAxNZ98QZ7QLzt/jtgIz+t6rfzIM7pSDKPhI2l4
PQJW4rkVczdbiApS9HrsS6OVh6t2MN6VOd2dEUo19L7/1Tr4MQoOxn/RJmJJDKXJUqoogfey+vBJ
fbFek88ACsyZzEKhpqQlXve1HhtzbyXbilIFgSuYGwpVmwY4F5Av6nzT+EYqocFnDOTWsmr4rVIz
7pPk6j+F/rIk/RnFCXeB50QCp8X4Egze/0kkjwD4FAUoHOSteFUuYddO5TIHK9PLVFTtnbqzoH1F
7W1r81D3r26ERHGlMBte86FYmiJUrl3jEeVZKXYFzj1mduxEoq7eAhMG2v3jr/dMerAwq6IOGbG6
BwNMSdGnxzXzswcs/cboJRNplqLS6aswYBF+Z+rvXWCXX9Cgbd+ID5b3ADkFiAH/KSqfb6cdLzTZ
a9QpMzhOfdHEH4f74YANvQPe3j+WjR7z8DbD0ToCazCeOnCaVxuMYegMO4vYpKAepeFEkW3xss5K
DCi0wANccof+WmA06m77k30r0h0skejgSFa859/LzDsqAtit/VL+CP7RZG+CelrOmSj+2ztk9yUu
lybQUVhSe92tGTZzcTley1j5C+kOv+FwlZrheijBfbaJ5teFVsnMjAd6oZ3QMYHKK13qwnfVsCat
M4L0Q4AYe1p6ot+UJxhITe8PXJd8rSCzUTYitWS17Sb3Re5hcF4whzmuAEgxYWrkzRh/1HchIze0
V2nKtpRFg/cD1dpsia4rWgVNl3O5JQQgHtHbUfpa8NtRsLA8kTN6cOPFkO8a8HsZAdWRLf2sYqv3
LweBJI67ugFzL/xDAxY9oFBJ43vkHM3jn9L7OZNKg4p7tfgOy+SMq/qFUwwtbEjhrUuaJEpLT/1J
KjRKwVxQ0tOZxZKkwHwUOx/AsnRa2EYAjfpEhasOHuj2FyzkJpXSzeBKxZ3hBduLrPRibc33jXr5
8PbWrdYCjiyGl+6tNV3CqDfs1JJ8dlFmoQyqag7NQO7gb+wRhu+MVo7Iv9D9VIY82K/IQP9CQzWx
wsVDKecO69s0i/Yi2ACvD9ClF+lRVYvhSBAHCMeYCoN0AkuiCtCjD6z5Nv+jeTd3b2ACRlbiD69s
wfja6uqcUj3FFztkR4k3tVOmWVNbRvgb3jtvHUMiIbKa48AoYnC9vUecQRIL+kp7KA4UKTYgM9rZ
g354EYr2pSUwGab84ciG31HWUxYmMr7jX2nNG4ZYCsSZRv5eqKcdT0bEegorUyCPTpvZx/yzaI2C
zMs1IV8myI0X09QgARnbytpwjnfNR16bc6k6+37cQ4CQMXlReKPp/nxWgFK5mi2Ece0UmbMPO6VB
TN1jHwBcaqY4HcB0Whl45pbCua0ysK9rtJxkhm6t9cK1Bdk019549HDBZeXz6W6tpnFzhnnkiqjV
FChlcAugxsPQgpcvOYD7dh0qOlk+ioLecDakERCuK58lNfTfYnvt1adWNyFB4mrvobl6mHjuteVg
uRHA5gcNRRbcHCoQso5NiA3z2LlOOpxiOBLfuW4bEQ2YVMvQ5KOi6+7txZEvGQhvDwxskgcTXvZP
icSpzEvzaqsTfiwiUaPFx1F+SNMSx+Qcajl2mksolNviJHNxwGVF1kXCRJUCE36+UZ54ju4Lx/IQ
eMal6oUfv37PW3usgmD8Dpo/XqhsVG0otrTOwn91dRYtieL+QtlzeTWfm0OQUGvrUQVTcpTckNu1
yaP+hp3i0huWSamFXQmqjheV2aBayAtRcJSxRoX3RxaT5ypKDRNDxavH927YWOmPklnUXjHk62jb
3m6D4y0KcTIFVRUrSRz3qJk/tLt5IrHk0s5+QUMX/DQWabwo+7oxJ8egk2ql77Od1/ax5flGmDgK
dNPVnZjgRNvVD20T+mmAwfKZCk3R+QuW6mef42nlgNb26TLfuWj0chqoo9yg/qqRxVwPbvtJuSuj
rE3OrQf14lV8Vx5SWhMwTTaXnJPfZ8nFXvI/Uhe8Y6lBUkFNye+Y40ylIcbcVJWjuEXT9ZfWVNWM
fXOslDHiKfZJ/iACQM8G8rjS+I8biS58rbVwksb9sBmMunGJk2k3i8q8bIWkXdkgbxXMHLIyxMWr
I49avUdTw11cDqEpjG9fj99O1VdGzerbUKyHiukGHZ5RoyE2SG5ygsqFIhjyYZ7ydiixNfT/9VJ0
blGicRDixNDcOg/WPqjUlwOzTQJO9wKmhRLdwrYTf0VArtl5jXuDypEfkrSdnmGtykJsyKelSJbk
DcqWTvScTN5/rAD6pwCAaySQtlSvZcUqI1DQ5reu1D1DqhkobgSaGPft/NeT3m0wV5/3JfWgSjJh
6FEjl27LLDe6Gzu/CKEHH9NM1mcMK09vaChTGFIRCTStU1wzLOIMUkHbaujjWSSNiHkyQ+jYaLuE
UTQngyZ+mgmL5aMFoAjZyNEi+N9MZiaCjEjNR6pSbGmCfzEVXV7IE+bFz1ytqCAAV0dBf1FUGew+
F2Axqkv5yEWWIA4Q9ZwABY0EpQaAJLm6r4dh4Oq06Ed92EIQlWZfXG1/4zH51ReXeWyNGxUyfsMg
WWOHupIqLWORX0kHooByAUEpnP5RiPC63uJzMBztAVwL8rucA7ET/FbpuMefk4qpw9oqpM99lI6X
65sEfWJfBdyps21siqrozVt5GjddLqF3BMWlpS+fyAoWcjvFPWuWjbMG28tMX7k9Vk4GiD+sHFxY
Xx/DBES3m+hrDDIlujQVKBkFd0TXA1PG4WyeKvHNss07Cv4zqMIviaNocrog9tO0oNtXInRVnROh
3tbcJK+Td4ynClJtLAOx04lyoj9yClYGNAleHXio+fZiUXLKIQW5zMSD48XrAvY0HUnGI5Avge6p
ZHS7S+eDVWJVUPaBtNDHPx3YR1pUiqXtYYtU1V2h37lKHE4CwiJrDzOiO8dDGhN4o6xtDWtjvalN
CP7tQqK/ywV3DsHVoG1WsV/IkIG+5HHSFjFdcXjcJNC08xsYbTwaPiEWSgf8kV3wK99SGh4MIyIT
yR2W/hWrDMR0D7N9M5E8vD82ZTTO8uMCOsimjKs6qExUuxMm+ziR/yF+Al2mjobAx4kuJQNErN5p
4g+vAehKnlRsIY2ksvx+AVaXE5c77w4rJAzoqfyvOlw/zMxxD+hLZLqkR1iG9fZtTr9XVWGrYsn3
YrOEcoUubP23FiXMbqgc57kSQH7NgFY2p5/tktrqZnFBr4EsgCnvp8fsMinkpR1pgvPtdxOUQN1d
aV0q4ALBX5KTc+PmMC2ow1KimnBE5cCwqhNomNg9NIRs3b2A2r36cYI52cL3nTNyZq23Bqk7/pta
TweNdroHY0raCS26hsRdtFLN3D0JhJZxyoSCGBQ/6Fqbf2XMGLeBP6gtXNd36vbJuOSrFz+cCbAo
EO54nl0N0mHcYUTu98j5mpHPfLi1gKqnb2APHIhHZBwrca6X0KoBq7WW2BXwh+b+zuf7rMCCNiy6
wXyo5Vy3Hapgf1/LA5wIdhbyVIj/tmFv92ZdEB8NrYHr6vJ3k8sNZaqbfUh0XgL9Y41j7eRjriGu
2HYlgK4GxTGm1tvwrRZxZ7T83CZgVvD2RH1O/aN4PI8j6jnLacjKOC1tKk978ikNuGBKthT/8cFg
clCSmcH+gm+HZhXcGpmERXiE7a/QTe3RLWg2ZkG9qZvrmO4trNnA2zIaxZKzBoJ8YfSTFZAF2rfP
XQ+0tnj5lNZZP+1OnugbazXHRIEwdunHSzgDKYUkrVp3YVVWfQuq8iia/eD5Vj/2L72zh3MYNHat
zS2OxEHkjdxqshbcrJWTc/zGfasONdDSQIxetx2NL+t55a+TgnidMP7nhU9UeqzoUWfThDx0wwsJ
aBoSV7vHa9y7RVFPKsAzVmId57Bjw4CLuKDRuEypeyK1ZAAkbarqMLtFSgmugqqd+utWNTdp4azP
yrFnYRibzPMCn/oI292Zptkkudl6g4Nwi3kkpUwAfcj7KWAS3NQ7qkx6/3WlvvBOAl/r8qN1OW7P
Nou7017xE0RkkZeRwJWa6vLUA9LVAmTc5GjMGurxrS7POh1kkbh3hKHZH5leSj1O2zfBD5TUT5wD
bfcecnrsucMg3iUBdKo7JhC6zzRRCEhyQTFAACKsjoV779xMKWlUjRVHikJkeBfqLMTR6G907lMA
EcqLVKUVTQSfMYL7Wn/wABu42Upv0e80MtTQ7l3lE0MnsP82acgIQMjKEH31IWPWURWgyJ9Ea5g6
r2R4+P8FsiokjZlU46rp+udB1WdQRmjmvuIP3v4HTgtdurmo3scoMRCCdWOzSdM8aXgdBQUO44Ph
1UOubO2gjZFSNAQI38JN2zblSZiOurw5OgSdTQuNSqzeNTwbLC0XuVTLRPix+vKHi+7yIH6OGFFX
j+6ldhgb/FmO+TU3xdltlZAgTi16ZBgt5eluAPL09wguhOlGxfWPNYFcAadiy2Ls3TKeFT1987UN
TjnZpp21b8LESvbkm/zGmRYLel/HPyTZny3czS/OHMsDFPpzNHqM3ofEjXOdWcQxROaweFM8dD7y
yzarqGYKY/xW89+3fZA+wnzkyDYIGYDDtpWF6aUme6J2j5IbNX4dje0WXQVKW3Aac6rgGfwueEZS
q1e53ywS9t+Iv3zF5wdp5Iv8vyVkq/eVxx4lEDB4wzWf7sGacjWxP1cHQk74V4rLXaifQqeBf71U
KoSJuaG7pUCqYjkdieDlsscyY1PD1p52VG49UadX2n1efcn67JnhA3K9yhy+Pz+1zV9T8UnIDsLJ
61O3xhg6X6UO8ud+7VRTvw21I5eOtVavkxRfCvtgfOk13P40V8X9IvOlAsO4jTyqzvagc8p35jDl
6gc+Xv1gf3Xw9bVtayZ+KCscnMRmCImT/BzrQgkr17fUEOPh6BgHBYRFvyCSIMcjupAHlf4PgR6Z
DytJr38b6TRK+nPgX/A0yAkOkSGguZ3n1I4sTn5SJunWF317aD2CIg6kzqTtzFOYNlqDRfNF0GZg
JfHIMq1DQBvnuSmu+cZN9gyMr7jK8SF9ELlmYdej2bmgYozbLdKmBQwuggRuLKqcpicuZ7wYlcIr
u9IrPFGGGVRmPFKV4Mn0SbRJjSa/XSUDo9CFLw5fUc2/NbD+G5qkx/jZNe+rgif/w4nJqaU7I3Db
JGdf4q9/Xo6dvLpM4jEHKeEhYefmiLQZB/yrRsWxLUl2C8DnjFOAicg2X/wJ1KPbJ9p4mlW8yy2m
rex2kDAtZcZ3rYj0ZkEAHI5Kan49PN+pTc+13q5L0Kn5ZeuHYUm+3/tMaBNcelQfehJ5SpQRMqF/
RUT+rlUnXAMyywpU7blNjFwyF+8QJSGb0H050ztZ7834X6ZRAQwF4i6gjgV8+q1Lw6ZUAF+EzPT6
jxAcAZQD0JjQODre+6NCxJppBuiZfODIKPxBgS6s5ohrPwwUw9Eivuh2+b2g3AU0ZCxRIkIdFfZu
LnJe2+SptKlnArlZAYd2vpx4+uL/knvXRNtjG0ZsAt2UflBXtKBL1h/xjSSjQwFfL52kKE2y6nNm
qHfuhxOswlidfAjRsAWcRI36WJ9kNxxMlxZ9uYsyMMtGJ/N4yn70BKooCl2EFTwYUmSVYzc/YSa1
4AldqeHQcpDU/SADcxS1tevCEuCjc3cQx1Dy4R5HIyCUsYrwaCh8icoqrJ3JgFMSzJ46ZT9tsh+C
tHVySQfJ8Mlj98FphGePaupSLIrtqFyDjhDarPejt/J7cj60cGaS2zEmPARI9xhz6nTCWWuPPPNa
e78PylOKajWRGBU6VIY/or6iXRRfkoIPShaSSXAbr13ouElyj8uE4M1iyQl6vZnrfiX1v1FX4GcO
6di6GBEumDHVlKRZkAUqgj8BwEqhAXG2JaszoiLz6mz6NTBj+bm/rwhClJjh0AjeVBeUN/B3R6F9
z+rKzl9j2frAscoKK8PaJhSSvWaoFyogWYZzu5vqoub0X9bx7pMySQjQ50YoT1W7OPuyA8U5AphN
Ykh2YqxALWf6rM8TTPEpBUVbHyHSKfufQF4q3ZB4iUIn/6zpxHMdoLTmglH9H/0zj63HBqB3HAnw
K4T3di37kxy+H2IjkX1X/+Kh1E585rJjy6rpnepjLqFQ5FoPwgL3oNu5uT7aZyhgQ8LFET+mFu42
tdnSzBlNEr//c1PAYJZKDXvkpm/7i5Uh9sUkjc9XVSbUTQahBJnW4KV0A3YSQPM2BGT02gGP2bdR
uGcB1fcWqUx33hcgTVyJViSE/ryoKHH++N/B3MWLehJMwZySCt2bot90yzhoxnSmB53VcDzFt31x
3dGObxIHgW6mXQm0zTkdS5CRnTlEvj6kTRdZ4yGMH7/FHtRg4RwLoTMdtg9+K21q2B3tjBohsjX3
GTmuhdcm5ne7t2aer/qhPi/ymVWEkaYTmJqINBGlzDAL84c92Me3dY5lGHOqxrDNrsdXLS80gskD
JoiTQt9lLN/BmBo4L0P2Kvgkl76gEU7sfzm5GVypIyO58b5ngpLWQaksplwhkwvz3CZnvRlgimmU
7hQHtm26Pu8D0/SkNEJW/vBUD5NdkmY3IlOW9GJDlmFYSnQyI9uifKtjLNZbz5wIwXun+glNKv83
d3xuQfu4nlNhgcV4oCYTxwNWEpmRYxEhKd9Dw5y7mjUPDzhDKu2HdWKH9Bj22G5uDb7euTKLeVsC
wWkGJQfEP+LJNerIwZOA1WV3aYWI50QekYmLhv7XhIbtyjgiIBR73tQxErH1Ib8aWLdRCIMDBGqr
VHJYITFhazc4xLTnTmMHhNVv+Swm5+frxgfsBTwNTEkpQZeL5NpxTDx+jNAg7ALy8TimrJiDe8V9
x1S4z+dMSidQ5v4gj0+ayC5sIexlq0IJkZqO7AnNGQAIhhIQuT+Fv0tT9j7yx5St3RIiKUWJ5+mY
QQobsXzqFCfWOsP5d5UyUY43t3BDm8GaUjw9s9K6wVMzyuRYgqvPBYs3ECZ5dehyzR7xmFo/kmhU
+WyvmuOinSXz2WhH1uuaQmCH4iyuzpG7QC8UfFO/QxIWfDD+XfQqaPjnFPBLpiCzo7nWMsW9huAt
lnFxVpl4mh+qnzeKS/tMqc85I1k6w/VjE3dfgBRtTUMKuB7Pdi/EsyaEXoIeSw42XnSINgbMBeGn
1BwYjdGE/Hd8yc2bxDmUxzeQtnxlDD7FBL39w/MrbCpCDeYAGl+unWoIzNzW7FZLtGOU0PhqlH/c
cy7NajP+JFL633ERrBOM0iKwoYr2Tu9uHqEZgWV2pc6KN4ViZXL966QO1vg4uJg4TTQNIfv8ZEUP
Xeg6lIhDkICcUZBNtIjwPZP5R7ic1/2z/wm3spv5NDq3+J5VrMrJLMC1a9pLFNSpDL15DjxLY+2h
3jB8qtOssoVKRjdqVkoGzV63tKu4wheAlQ2Y4zNEwNsjJhf5qPVFaZpG8StjnE+VixWcbP3nw9At
PsxzoAIhoaL1s32i8T2yUuVVJXGy3jdjCb3cwRGzktWvMr1sjaHpkY9VFyOphGL9AEVZmxI+l1mh
VT5U5lLiOpK9DAJprxLziEHc4LEf6o8l7+qdEPBF+TR/1Y8hHquF/zU8z9yRJXxIZTTvpmWznsOI
/PPBvy8bXsUKBteQi/EqKUeC71LN4ebgUiEy8V0euOp1bOLlk6Lqa/fGUjv5kgAhIMLwtNeQP8ez
k1bCY0qNDdrT3qNxkycHjKt5kYHEiLMwR0ymU/DFhD5OUeK8EW9MzYt68h42vHca1iYT7uYMXmbM
fZzwNSfikjc2y6cpBJzftM6a1eFr5AwJiE0Utd+TTqVCyKIHX7EQqyZuHPzxW7+8Wee5ujgm268t
+ZkPkxAcyy2Fi9g1J8mwC5fZZfjgJMwoVPVWkBCYSGNyPeSOA+yplINWx9rTIzKrWbsr3lw4Egpq
MV7WzZ2fUY7g0RTlnXm/v5T1Ym/NETXBeWTTcSYxDi6jOo5LiRoe3hiRD78v+OwZFENPBfVX8Tmw
jSmib64MG73mh4i8U9nk3mHUlrYw26S5GLGXtD75tqsPOvSioWdt7orkDvkM8LnP1T3eeIlqGz6a
QbgruuZ/UghSWoh3ENCj7ZOloQhKdQXpKaZ03OHmY5adRfD1WXyffDB4R/8oOwuTuLhYnpQopGd2
FFNxN1Nokl4z/JwmOkqDBpVpoTjEbMYU//6Rehruv070LxTAlvBpITpem0NsgSSldINVw/cn6A7H
PFRT5/8gDTH5UZOQgRK7TDTRp5GL86Qb1Ks6h+p1UdsDayp7c76AXQLG3HeQdILhx7FY4Sw+Pygn
DDWQQkb8hRPbmBwshjREG+hnNFnqwi77qT4uSG5pIgZnL5fcBro2PLiYYv2iw+2OaBpviQj7PVVD
rptSJAxYTZrQAqd61uO83hstd2aIY8KlIkkTISHOmg5Se6W7trorSPW140HufLu3VGvgmbITu/q0
F6NdEc8maGVEUZNB2qRNd+YMFcX4GQfAJP3XAJe3eyyyVf8RUxzhmPGOu0mEgFrHMB2mp+SxlUJE
TT2hcC5NbFL4hpdn//NrhavCmwfGpMd0l+FYb9svx+wGsElxlEPm0pxH/LmPB/WdU6A361yBOeAV
vt4B23RgqqAiG3qzc2ASzyWR1AbFglhFGkTTW1ngGi5W0EtHjzAOKZonUg8Ad5zIMIUmvgYqLYyH
YsGJuVRnVz88gTGr9jPi4J5+De0CfrsBwqYTGZAaR4+InO9ta4wUrTaosG9otGNtgtgFreaHscvs
vDViK7kYVkDu4VDkByOUfTJH6kz/UsdM5hk8kz/US3FBw9cn9ZqdURda6PZ93Ldus3rH2c9vjOIw
ONCihHxK4OdTuINCjEkcZ4Jad2rg3xIrusQ1QKW9fUdurQSUilfkTEn/V7cf86Zt453kVf2ZfqUC
ZKnAvQDPP9vgF683IF5QtFokmiqotk83HdhfYzkSUYyAXTzkiwqz1Ebyhd0fuz/fcV9vI0aOaBJQ
rr4J7Bo741esCmkuP+sGbqsfWhm56nwHSd2mJhQpe01atAnxdz54jWXnehymlbGVe14ggVE2c4mV
SdFWcVC6hO3yIoDxetEtuA4ft2hZ+quT/WRJlxy2eijroxlkK3zLfYXcLVX2rd/lb9EyWfZDtEtg
bIOCc4fREftbEy1C/3wDnafvECI//zIPtRTNCE9ht6M/AO9cNITuEb6YMDmAmZ1dtUmeHI6QXlAr
MsANnxaEkYupN6SUReFFwr6WeKcrG0X4gtn3weBQB3piDm41xwkCJhkQOBt9Wk8A2qdmdH/u1us9
ffd2QONm1MIs5qXki43rLYjxBbMER16KUVoiMtaSdr1LL+CursHgHKtn8xgpavJXrJjI0JQuPQQM
Bec4B+hAnCo9xp3wKMi4Kq5BJT5Oa3+fl4/sT/ZUx7gNnmRJQynbhEcf9CRcEO7sE/t6+0o8CXti
odO3FnSY8Ubslw0HnzfWZ8KjtSFM0dquJAc/Nz6Zm9uq/jqu/ghLYgvt7shIG+3EXtz/etkWOcws
TP75RHer3Qg3L55AaxUpn1yHVZWyEX0hlhUk4k1lTc9CQ4I0EfHnhteLdRTfHdrA8xFgUjlOvGB0
wqoDktv1ioPm5KrID6TtcxiDFj0RmDT73B5KJZKCpaEC6+IPxkoCuKf+M2VAX2gBhRLDExvCDb9X
JpK68pYQLtgmxmoJud1+/awE80j7FKxIFwyggLcBeDwSNnXZRhthv6ps8AKUY8wieuWvomdzYr16
4LzViDsOmxipZ2cBALFSpGC6jgegorYRJMB2AbPoniST1zbl0YQRILd9x3qr5okcyOIDF3B/Ff0Q
SGT8RzLiZRk8piQwNC26kJb69zAbRkNwXo01Q1ozdeQj4rV1RE0MZPpbky8CK+707FNKIhbOGhWL
G2AiZRt6RNDYWqDMJpwjE96Ganc5iByXPhvEU3pVaimnJXzkwCb7oMokU5GWYrzQ9FBAfjjdf1j3
L2JNLla1JunoJMJMvhdlp8Nz9HF6vPtVzKC67CmqS4p2DwcMToKfG6dSl2b6dQZJD3hjd1wuSejC
TNQ4dybkEVyYHF4f8F7SzthlpDHCmc+GFfd8oqFFn6d4+pAm+s3c2YNHZzpqlO5fpnNPFuNtoWef
haFhxyiN9ip7ZVdxs/0z6m/RGNDzDcl4zppNBN2ei7RBemTnnmtPWg0d0e6NuzmnBSiDC2ltORCp
isHHR1aWAX2Ja8D32VzYEyyE5AMk22OM4LwZePXLK1KelztYSXI6Qk67YDJz3VsIurAKBVVJeU8K
dhOSmwX6G0E4K5+kAf8l+ko8DMViOtDsxqwgD8gQ3dHNCM5PNRGj0NNCEpsMsVTkdvOMn5QS6sP6
oKyyHYFDZxEIb7o3XwRdcpDcaHI2tDhCABhWAvh47rD1MZIGbS6+Aip8IjrE+GFWAz83MquC4alp
8w6jkcs2gJ1ZUFnVJTEcaRcyGXCM0DzjQSeM9kFN+d0JkfA3uDRR3VuEs5Z3HdskEWgCPFY30FOM
ulXHM+wYoFV/kdDvIAVWk+W9eqEDk2Y4i5Kizaxz2DtSVLf0Nt5HQfxcTbGBm9YXJMMZSGBAUGk8
MXWP/ecY3aj/9evk5zFTsb/yPWD2OTg3hnKiTzwxe3Qbo91R6/BC2k4TBVcFDp25wKbgLAnulY5s
a/4fA3DUO8ezsQgcfjm9qMW22jL3+mOapvToc84PYz3uZkBd8TzJujLGrKnzahBglgxK//CH8Kan
MSaT93BM9pZE5b3F9q6NQFkPQHJqWJjhlidB4K8umZUmo2hZ7NpziTQfILUws0v6yyeVzfciNpi5
AwW6NNGdsCD2xNNH4FGYGpdYex25e9LmVq2DGsFHaRkx4KUWOT28zuhWtBs+1J7n3LkyFr5YbyBH
8Uhzcvw4pR1hQ331Xrytxy0FlqMc8Ek7f8BvMstJXmwrWp8fDnTWuKKlDkKJX1kwCDXW+24WxSF4
gXPVKnP2R99mT+VkPKny6YEFLmzNWPdPU9Tz/5A0ZLJUIfH0KZhhzuGpauwsY8UR9ihKsZLvgUg2
cD0OocMWE4/Mbo+iaD8d57ZALWCF9xAN37I15wcSy74Cfaqp3DkINeXSlDYkflbtn/ZYtU1ERzMt
CG30A5AiOLUBJLUjsvLhyMUhHTG4ZRUn4PmNrqX488AL58/0i7xmf87gztB4wPPB5irPH9ntE6FT
9y1H+1opuDuxgGbGeCG17pUML5P25eF9ah9ackIOs75YxdSLxVsZ9cYVZIeTU3tXgDZvNLCHL81Z
dltoP/kXmCc9+zSmqEUnDliX96TokcpRym58vdOoj8EzU1YfPxDIHkwsSoqFjCAvs5I/7lVLAAib
+XFLXXX/EVdJUFVXdUZhpB/mwWk+aeMvCUhIDArifIfGTW5/bN+0y+5SFKVf7wwXZs5Yia32sTNB
xKOeMwUjR5hVlNvgBGTarPSlmiT6UyOR654J9e7Zpc3kSyWmEtCn3a7TkxT1mFYmvhpyuTgyjWY3
ZGdhd+9Z4ScCQVEDc+ryoLC/W+YBLqKNkkSIuDAePe03bFf+76ldwZz6oOMvWqQu2xq2ktynTSTi
xaUnKUkYPQlhIKZFv4qpZZ/6NRevV/tsdmf/g94i5cw7JBkAeKV7SZPG81v02TeyS0hsgX1AJVOM
RzJ9v2IP9URC3B1Ar+Qe1KSHfKAsjK7FBkxYPiut9A1MjXL5RQ4+SbMfBXr24GHKCCGFBwmGx2Y4
uL1s9K8AjIbs+DNf0arF4g1aYixKmuQyhfUw0vffLXz0BGEpr3FLhG9cEv2qrqsxQzSxbKwYW88/
Qdb3qO8Ko3wO8kjunrVGwrsaTm0WBRSXbLQOHXhygdk0kdvUDRsKOT2bPWE7fyQxYEyQVuX9MrGQ
o+MxXdrNTsOBD5Z++fsbh+83xQLo2hyFsyI0u8lDNE4vRYfWFfN+VehMEUzi2kGtrzmHIQ/FZl+K
Q0fi23/xixWdaF72+3sP3GNoA3Sf7B59NENP5FJu5Absa+WSM4iBB0N3mefhLrx1MmByYxxAfuyO
luq3ngw9QK9nrQu8tLk/Mkc5DlQ8zLvCTtiDw5RxXp0hlu3dTVQ7Y+vhZx2BjPruRvlU2pNaYdQB
W84I/Ylss8mb+czXSlGKIUTX6wBbIPY6h5dG5WdRPYVQYYP+xu/r+qhOvdqkIIifER+EFzHgSEMB
3B2RSer10xkb7QHtNwtaH2YM4vtddLJGY9Y6v/2711uwdsdWIDV+xonhsRX/ejF1IMDnEDUXlkeS
OpWpuS/PleXgNLT8xaHVHczMI55S3Za8nsmGenEKmH3xJTj1WCARy7Ksv0mDb5ZYFxtrGrz5O68n
3nYWGtZvSwZja34aqBHB54wziNy60P3i+Dmj+weqqUZl4rL0BINJG/5MPMlqV17eeROFlxdyutMt
v/5ZS5n9Ot1UICotYhhe5RL1MaSSYVWmiiRhPzAuLv7arZI8+ueSN4SK3QlEI+f/AcFl3OBcPqEM
AkhWuJWo8rHbFMZzGhLbvHk/rf2b4yg+KPS7WQO4w39IWWoq6jf3r+R4niDBz0qE9d5mMrBLbPhx
B3mX6kxskgCPooJTFXi4wDxR+HpM+9OWPSXdGw/FXmcOxYC3ia9/ed15FF2MM6KNb1ElyEZqgggx
ZOOnCdPIMZEp9RgSaATvl8kQPzskEy2VhkuWPTD3TvhSgY/slf38xmbUP01udV5GBeE2Oob2nSNQ
2c0L4TYJz50ByCbsIXEbM6TJc+zSlGhaiTQorjtRLTfsdIjo01RFkuifel7cHYxG9LCKNlhoC3Ya
NtbyR/q6fs163deM5YPOmjhbsqxCkNPDWbzXt67zNxfAOWe9B6i1BqSkH/sTptQ04WKWZUXp7FCo
84dGS036uXzn0wlKj780lZz6Kr/yxs+F8uPA6i1533s2KDXrFuNkBJQRs1gUy1m+ZI9St2sW0xD/
V5z6OLR3RuJys2MIKumqvS1LeQQlkyAkWu2Pp9X4czeisGHIZJ7vaKk5eIBFqascBkywn5Vcf3sQ
5axKcOb/Pam9eU0NROHOGeD7U/WI2CTv2UEClXjUMFFrZVa/kkWkXf/tm/wiLFvfV6C6vS23oYhq
zfo31uaLd5J2nMx5Ftmlu9TYR0W6RoaJnVanzwM+8oD/9O9MmenDua0AlppjiaapDYW54OdoRVSy
GlLVETbzy3RkT2P85SGa/GMkyupq71tO6ghsQsh77kjPSrA7a3X69lMHlXnguRIAqOTkvTQWtbQK
aD1r7HxtoiuUSqtLWwxb66ouoGRxrl7sEbwN1XfrQFXt58KPy567GybCYAp86HKz6NI6TiLCLyWh
Hfhx3P7WmjIhAHCD9dnZKYX60eiEvMZYTJhRLk711lXsDvUXyOqgPLgB/t8ndnJ4FsXsUy25C/5f
6wAlWL1yXTh/xB8VsnR8cnqaBNdKs0agtbedgL/3ZWv+EDDv0nAuPuh3itgoYjmqdu6aUjm6nsYy
uZt97zngrt0EOOjDlDMGX1aLxDEyJVV0Nt0BMNSMaVyTSdEXM29Iv+YRVRG3GotJbgRIPs2g/I+T
a8B6YX3c80H5ZCIXIOqj3U7FEt5nouaBwmy+g7JeT6rNrW7V/7FGybyNXjjYx/pzK0+3ygeaN/GV
+zTF3OnoXqQSm6yfvFZRtX0SQ6Tm0Ap3BxzSCRFfJEEow+TIbdWiihcjR4ZtX6LBC0KLoaf6JFzp
Kn/6+C5L/wbnjKJegXmgZTcPvgbSY9yBvNdRYFf3+VXvcB7R7IjMKkdZHPyCTDbyBzXGDayzI05z
M3Y+bpWrNP7epBDGkheYy/StFo0w6JtG0aII0t+qV5/ML/GPLJ5U0SJRmYUCpNBWO3PHpLgscZRQ
cBaRE+q+q/wTvNy8H+H/wRbyQLY0xk9J/gmp6XJjDHDS8F4++x9gQ4FH4TX8HSUbtq3SIBUJaWrl
lx1k6tbRLCuI2VHgfF5LLQ9WAis30hWCwQIF58TQDIMardDzYGx8H77Sj7Lk/qBUXxEiNnzH+nED
KZ0v63WcPO0jSIl9iBmzzjqSWPfdHFHWMwzWL3d6uBW2W/yQZXxhM6HSw8HzAJMkkMrsKiBhIgrH
WIBQCdK3xmh7sHKCRq1xZxApUaqSPspwx9MDSvJJhTBzMZY8+/jSFHHxnSHf52rQ6bYKpuOnjvRk
Zc/uw1fkxyDSmLlKMVXjCkU52ncf2iJxiuyeVEg7pkHl5wWtaqXKbS15PBqDqCZjRyrg4pfZ9klN
YKSCEsKPd0wlcRKTSYzCFao/xrhtLga6CChWX3XRLlQMOfOiBaXkpA1z7p3Jxx/P78U7tQ5H3pdm
T/LpMW/7ScUg+T4N8B1K25fszlgonL+PttCblhJ6bYGY+5S1vRGFX7lJhXNb9NLjVag38Kqpl8rF
800GdZruVq/qrOUg66RogYTMCrkWY/9H7RIpsanIlR36PZXc7TBQCwKfsfRkOpKM/mlAOSz6fhne
K4oNqlK7xWBq90CN1BZunrUvfmCXBozHp2ANfDXIT76iQlQciFFBgRV9zN6lkQIc9Q5m6KWEIzKz
053TstRP3i8qpquje5u/PeyhnhWkN129ygYalht8fNeawckzyPAzr2hNfM6Y5/bOrPzKiAvPDxOZ
kg7GcoFhMa1IzQFIUTLHQf9Ugu0feKjL8Arsgdk9AwAEBo/Ue/zdQBCdZ0g4U9N0xcbqNSoey86g
rx1aH7eoIC1AQiLeIj1QsMI2jTewrHLLuDtbl8icrwT/nHfyeONXx9R+7uztPL1c2K76ID5zY6+V
H0dFAw6NcQP74GLtyB6x4PW4DD8jzRPreIpfyoRiYiJMJPGn+4fOEPXpeOzrD4QMQd6WXDD/SiA4
2P2F0V9Qr9YRtwg7tSMIcr9+zlgGSb6prLZKgXUVNl3Ao3AfX+Bo6jO9ecac6D1VgKGlYL6iX4Kw
1WxFHLOWxJiBGxIPPToBDRlcRV+P1e2NklLJrqO/bTMZg7naZalHXdLABi+QaVFDphjlzMxKhRdS
Ahen+hIvHXKVgqWuQvycpN85/sbgVQJK/qIFbxXwwQc1pS+2jw36+Wg2jnxHKxv7360+V7u/8RoJ
tG7NDWXR24+TH/qrFztn1mV2XsbEPk6MbqsIJ7p65Qcj7XeWRpNxgT7BIQ43hmJy4Lc0C2nBXc8l
TD+UeRxzvzneRPu5ctqiai/O87rnOJhe0J6Ptibrbgm0x41whWKOjaPnrbuIVg6Nlpyi1OSqzYYs
D6AMYQSb6RBax18ievlX2o1LI/pItsLxf9i/W8ylgZUJn+LXYPxzv1x8v6ayJs35TH77hbZJvdlu
gLQwkT85o7T5urksKXZsqXXVdbGg1/hooUPQdr1CyOmaS+Hops3AnHJWpU31wmzlGw9DJPM128Fv
Q/WBklgW8JntQ5yxWmYduWYzq9eX/80T/2tYjI4YtKt2NQ9qPov/PLwkxsb4u56cZ7SdJLbVt0/q
DcBd4/wF7TLIwL0f4qLu8DmqYOgEaITDq/fb5v9k+bZhEJ5vXTPsEP/V9jPjyVMxkxGDGIZ658MZ
k4vQUeI5JugMlE28QAyfJWQXknDblNFUqRga/HJKDXcAs/doPfBPm6M4047AudtkdXLVbJkF6Wcq
PIpmj28GQhW6yUKWcMEGiicAZVEuZ5GUiBC1zjmoZVt1NT7he+6pFjP+DNWFbqsTIJezyV3gl8bt
4aqMq5b5haU58SLBUAnIcc7vBpLodSHrNIzgKkpTPnXKHvJ+UImfNhNCw73jrz6XnwYfhhf3R8rL
97KiV7oyeul5OvNxhgm/MDYKuRBNBoxTde6FzA2oQrJXusyVdjA4wrdG3LqcUxld2xMlK6IptriD
4gfNvmJFfZTQChDVVBa6OzIKG+8gQCKEzLWQ9qff00I4z0kIpv1AeyIgg795ivwrc3ucnSFe5Iye
IUGZPaf3l/+w2LXKkmKW47DrObR89Jq+upyThTxbuDrnHYlXvIjrtElz8+XNJBW8UZoi3P4ZkVZb
tR4gRUD8nNO62Dtsxa7bd1QXhsZzwT27FBFOiTThHjtpnA5qzV6s/DUuG0abrX+q4jWahxSqmSVO
8NlI0Q3+wMHrqsgGceWjGG/uUPmlM0fW0PNW8iDtIryrDerZQqq6kN5U7qCVJ4L+R4RuK/N4D17D
/VXNC5Toij4vNYrQtvbkFOI2rCqJ/IXWCJK3IpXXMVOiGT7Ajqj92O344PaKDxqsxAtA233EDXOJ
DaXgloB0igLkhwWGj8+B78R7+3UHUHDOulzM/dR7UZOqv2SG0Xkh0ggephu/ThtVlMN/PMZiyS5B
iHr98TLQlTzCa0K9CtvFoGLEzj08iCP1XuMEGYTe5eVu5Q+hZ5laJ7e1N6yGOQY6fghOEp+nJEKF
iRj3f38f8G7ZwaBVSgScHgOVchzWdBHvwlka1kCK3HmRd6EafUmsy0IagPtuYTwCeXOpCMVedceF
DSn4UMevFX6YeJ+czqZeqyqT6Y/mVnvQcwBxUSL2/t6DRmsK+6BxQ8Ji1dILSvwXotV01sQnHM51
/W95CS86TwzPLjmxBl/MSpxzsL6SGr2lVUjC2Lq7lhBrGqzepHJ5SaHOewsXI/7/6ArRRpvarWzw
vGaQDGZnZyGF8nWONV6RQL6EQKKmNXQ5ADq31OX/u+d9oHrXvErrCTT9Nv9TUJP9eBGwh0kdLs09
CYNp0v16N8UuNTC0j6MrX+K3kh7kctiW87mMezMeg7EWjlexQVhO4tumF0/Wzh0RYOgAPxae9OAA
tVANbiEYp5zunIs9nbltpYM1YJPEzAOFDmJD0iFzLOUqGwrt/C/tDo84wbvuXhcicg6QjaxgZmEM
2hK8t/dMqXHeb6DVe4+UsZj8Uui9AgeJ7lMlxlJpcg2L6oh0RH6qHDypjzkw752ovMPPXPbGMhDW
+6qdjNT9yVvDmlGWyhnSoEFMr1Ht3ytzdNHGcGS870heb2HCwxyA+z5WqxGFw7nY6GcHFrV1pDId
zE1SxoDuFX1OAx3ho33fo9rOmL7u4kyC/4Xrr2qOKzTkT+ECTJcc+xPnILHjzDCA2DDmBno7Geac
htaDTkdZ1BO2JTEnYv4fgU7gdMwTYpfO9A2QisjHKJYz69PSunLYnvkN7ShTbe+sigie21GMN3Tn
wehl5zYs6ov9tBy8ifl2JXcPncNd5mqMenByTpqIs1JbXEzRnMq8V1YekMgzv7+oAfVX9BfTaovm
wt4KiTwIp++QPD68Wii4XA4yA2rY7EOH5uYfrAyedLcvWHxVuP4pjGV1J1Tac6l2zq/6ReMlvxQx
k1xJsRp+eSVTUn0j2e1xReUDtV7wYpdNRfPro3TwvgYwOiPFl2VpU8Pt16yPGmno0zuLMhEawL7l
drmzYHA+B9RTzfsl+7WBAS4F9dtjTxRRaYiBiPnpaaYEmxdN+z7W0T8yOPDk5Ip1dOnL8vIgZxup
a4UiK8aGqsSg/fBjdnjvMV5xfh5/6xvoC5WOCOq2T09pqDneU2csApTDg33TxWjtfihkWQCx9GOk
tzsy7wEp1w66Wsb1yN2wPmg9Feiyk8NcZ3vum3eoxL91YDnONyWJy/AEP/9LYsqt6w6E3IiEKxVd
S3B5V0w7q7s713kw/IGMKk5YfdXibFlxk/lNOKbTm4zGIHBpuLpCQHNj7aP5Aez33+YXbqfWJGLN
bDMeEsiG1/DXh7QkSyThuF4wHMFJhg+vdK/CJjek7W/MMOFEFBM/cLd9ZBN8xbwKu6DCCFL//G7p
qoXwAYViF2M6wsY/WSrUum/IVP6j9r10W772G/1o0ZFdhbRNxjZ3jXeU9vzsnzN0IEWi9+eMLsKA
kgc2iGrGRP1UhfsjZ6bjfAytOoWp44ZZTf5zJPv+C6mWj3Eae5o0gGYw8pLUkD5ZPYP+iZCuQTPt
9HoEIH+RbX2I3By8N3JsZ0iidYZ+2nqmZ/bPJLMXDe1YiRt+6z9EdiwvQ6GA0Y4CMLQkDsBzbKiO
efywFyr2tQpPmJT9KF3v+CA7iVT1o3gEyjgEaVLrYvtUVgEzU60qnBtINrKmlvEIxSe0FIo20ilw
aOyZ/0MBVGlp9oCrSnxEc8FoEhGZXMnsMxXLKImBVhWdkhJSwb/gqptwnYkNPE/2+s3Wwg1uQGAF
z/JtKKnjCXLKlYu4Kr2arU+fDCtj7oj4jRQtkDzFj/+N7PfpkiW3gEuJJvwDRcas6YmSgz2fhuBI
nbjUUPF/zMWu6fljJI5lyuxisBZsjjSqTaWD1fBQrvgHQ6ytFxp7yBuByVcRuawvnm1ZFriD6u0i
+HTF/Qq5NkF9yyUFjpN6YnlS332PpAOb706ytvZH257ZDom1t+uqxT4+8aY7jTi/gy6zSIzyqFad
n+j7YpTXrid/WZmkHKLy0prFQUttqaj0/qS4ACQ0MgeAHPme2yU8NBZyScO1AqENSIHAu/YOIrl2
UDtrA3fmPlXcgb2QWZdsY2snM9HB8RsP9d1UmmpGxlwM6ggaeINOSnsL6lO5bq6moDX063S4cZXJ
OXmCHwGDyFQF0R/RyKzJioYXALCq9zrFlN2bTzZXrihMTZLH+8twXqQsjTiAV/MZLdMLtZllfT+u
+H5YbUUtmkMm6pJd9zM1vKYvq9EyerTC/NEYbKzuy/gpB5JRdsG8I7v4AaD+wUOXwPvamrVfXZSS
BGJbDUDvSSQjJ6+kWHQp3vLyAVzCiFE+iqvqMcrbd2zrI8g23IT6qCQJK5VnmeNcu916ngYsurcH
5n3Hb0g6HQZjkRth+7K1JoBPmVGCBf2qV3m3sbYBb2OiNqq44EJN73fQq9FlxA9SMxozAN26EeOs
jxxuBaqqhwCvMDZmyFR7f9WDUlMzhHcDphXt28vrfqSHlFhCVRBIU/Mg/bKlRAZSM6At2Eie2vHr
BcppFdt2zCBDI+k0Ok6VCys43/gYbc34AC+WXyT4a39wOztVFL5qGvTFl04JRjmRuYAvWRxohL+b
CLENXP7eZLeRbpN1y0ZL4H4/Ljmtxo9nBG74YNv3JiPgE3y5Qgaq8R5jCumGOf2aBPjfikkWN+7W
tbE6MUy04JT/3JxXgFSOAkC6S/J4zAK+nTE7qzUNDznco3wqE4Vu5TJ6ujKqhE6FrUAiUAyydFpr
pvvsThyFAuPCTImwYcCZLnGFpvrgIzu75v4LXsXlSWLDkvVZ9pBSCo8Vy3Sw10J9IONoAn4Vohfh
AVjyBHrYs1gXj8tGzkUNJ6ludWlJ6CZMoqSEnCqIECrIUcALF6HA8C6GmrxHKObrTpggvDdyRp3w
8s8+e83aUt9iP2Nu5edm9xeaYqCL1ds2pHZmENk2Muv19mzPcvdhztokuEq9cgOznkWKbbl3snYn
AfsMpWkqyFzo8RCcuLRwUxbnpMEf9fIQO8JB39HghBAbPypnvQVJ/xflljnRctuNJaes9SH2tjoi
v7kVjNelouvRMeDYGgnmT2vDHnQEf2V6omj3aJB+m0bQI8YwmXQtV5A0aUhjAjLNU6FDxrPofcfN
0PhvURe2pR6TL/NgKN1JrqyLQ3vAB3ueapdQ6JO5b9j+GCGuZzw5dhpxxGnwDZNs2a0mLPBynSLu
LPEt7o34liM1WMJytdJxqQ2q7ehnDfj09VczrQJ2d6JUOIBmSg1LkhyPukgHt2GubOg1mRqrUoCD
0gKYNaJIGqrwORQF6LgkRdJap0nRB713y/TwF49boXY1EI0/O9OLiDsSHkkJER98+uQ9wGQKWMeN
cyTjLc7xQYGTWfWZLLNvxp4ADtKyzhkO97iJhZnO5wGoH7OiCiOpOZV1AwjoN4BtBjgorOOA6q+0
Ln01MoPZu9Zs2NSzbHLn7i8FEAzXlgsM/20Vfa6op/REsWHweK8qWxeeNB79rfFAYWOpLRPEL0TG
ONa4LmNRslrWd9c+4MZar4Vm0LVpTg47J79Ill6I4QBLeHssB5ErUdZgO1PzQu7yJNcfbiyGwdzW
AOHqAUoBYKsayl85PRfJjUshQk52LVpkYekcd9LSRjr3kgqt5qqBRQ7qYTnyVWmfOxbE2PBwFto5
H3FjJ2OdBFey7t1+PTmw9BO+lLr7yloXAtD8m4P5rHO+GHEi/F1bYJummYqt3vlpliKIQKXE2tCf
9A7+X3DQnqhsPUJu4yhPgq1c1zCM9dx8oPGbUwOBvTTHdEI/3FVG66LaD5GdeMP2Wsh+GBBuH+q9
Y3EjK7fb7BODWO7gHqzxnGoZ2Vt/jVPOR2QO1cQ5RsRqmVamfRbj9JL7KnTz12MlUkT15CYsvoOY
rouWtgA2ScikEx6ZrZ9TPb5WEdSg7ohoaBegfn9PVuChWa67ChHPSYQ7KpaZDwNma3axjgMtjUyp
suqj+zjbGEMOmnxUx8stUmV0sHv+OQHYRURP64ixwcmpxfyzTGNHTI35OiUI5+CjDkuKb3By8pPv
gfZEERvUvExYnAEWlftpMeqjkncyX61gl/fSyTKSrH6s+/J2SWW/NMVjfszNETWZSQ4qaU/moZEj
5msWYVYKIz+5VB3kh5mc30ilkqGqYZ7yO7sSzwAx5XLv7jaxyAmgEGMgvksYrCPFEBm+z+OoHUII
FdjMpNgW0Vuqf6miZlFnhokN9qvlgGD+tTeks/7O4GvejqSlypzYLxzgv0tXD7Vtp17OJE+4IX6q
0yl6Y4XUb34a7e2Rg1hJ50bxm3rIaOvzmZuyELRk74w9CGeaPBqcwZ9h8me3GQFh7XUm1LUXELGp
J7QKBu8bisjDDB6uiQ03qfHGfEiEdLFvrTPZ+f4OPmNft8vicS+ysoT+LjIUkW9+6FFZF5uLUKtV
8AOy7b7zklov3/d8qcXi469iAjcB3+Il6p0nCUK36BDB2LLv/aRpEm4v2qanAPd5Ma6LQRBolESO
Bb6UchBziB8KbWPQ9OvIMXG8kxqBKr+le4G8As1q+tTHmS/+un3KfCzJkpCpjGF4W634UGZK8ub5
gofwZxL1+SgXLZ+pfilI5+xd/3NlmsLxiXUnL71cQMVJtiI2NcqsIyQ6JkZ933upwKINu4Ednbfr
wKLaMoZhsCbMjjIDP/P9nWYAyQCsZkHwqUiL7SsF+7DsGPBV69co+S0iez6W7o8O4dBHFtmjS5H2
zgE5rtxqFoXClqxLcVo4TT50Sii1gbPGyUwL/iCgM+V5t6y3z1jVLiHrS/+V3Uq4ia78TA6sPTws
PGFRZJSd7d4EHAEhor8u62zry/dQ15a9yvBfEAw7FJZCv7wzqtlhFVr4WJUlK7a9inm/DKpjpI7O
LOTIXESo0Nqet5YBl/nNINqThGBur+kHD2CbVX7/kjIksX2R+lul4dYxd720FO5jZlXvnQ+T2aSq
hgfT3UTQZRirV+gJy1T9TgALTyDN12uW2LXYjf+gI4Xr2lcDWXjTTmomIKj7aH0ADMpxRONVIflj
kH4iR7I+JUfaTZUiAbqUtywMa4oTeDxFA+jjp6enKSc1libpP4bPz+Lc6UbzGY/DRxmG7uiqUOMA
4N6A2+zO1qp6YPz60fuRYNP/Z/gzLl9j6QdYmUOjN/Ot9mJDERMKwzYwDriCgFaTYzHHOvF7E+b8
W+02cR7AdfgYn0n9VGMETJ3SczlHlvFM7qK2XW8Ntq7YR46jQ8Eg37Q1C4Vq8aQVvb7rY0LAuM8n
hVmQtDv3g1UWDlrQblmWrj8lQHmsqpeCdfwxf0h0qZXiosFfuBAbwnywp/PEK6jjgmi9znx37U3M
WIJgoEaCOoUoJsua1vm6B4NZIgQDHzDQUSx/BQYFG16qrjQkdD9m41GFFMFoecSb2NnzqOsAiqtm
hfGcASxQEYG9PId2gNlK6fnO7shhB07LyY/zDgorJfvCTxXixlBjAVft3ejrgxxyefOMIxlOlad1
BzaTYusMkBPbqth/AIzc0KlVV2YF5b9RN4u8Zzo8sV6Wg30g7+MXY64v4iFhq5ywoU2Iwdy3IWCp
eEzPABMsRawcuEuq98yHHyQ8dr0QjUGfJEt3PfU5dxqQ7bWrDottmiTZ129UDhq1JtV8gUgwruN4
HTlzaoHG04EJbW7VcjA/FV9e9xJp7WI7w51v831gjFyq/2vv8ePPXY37+A+QG+8SUIBXZHs8u1Cm
ua5lBPMrI/VIvliV7X0JeZ9G8xtmjsg4tq1eNqrpaQP/NJdkaXKh8kOUqWWW14qz8wN8Z6Nu9Haz
M+U9e2oIN/Lj4uyk382ptrYq2k5tr0n4OcBQ1j9DgkU3WFKrMAXjXt2+ULkVCkuTiF0XOo3HikVZ
AipArt2LQBenBIcz8sw9sayExoE6h+EU6nTWHe4ptp8Jj8c0Ek9+WazmuG6IRVlnTxv3SwMk4znH
rlPv8F7ARpl12fxCMIJQpAwY1I83afZ/xCDqQJHY0gUwgYisz9aCtWGn7E6hvAyrVmrzmkIQXCr/
VUKpqyDXpdohqKqnRQgA24P85DrQvVDn/7vryiO5NyyJ+9Vj1mDQ6ebaEJbTGzorjx5dUodmfd8E
TMUsvjzFNCW0jesFQoclbOS8cTaxEzRuVa4LRfzd1gybOLQqvQgmStltPy9dXxZqkVvBILTtugQG
h05e4hgLETlqJYmhVszAvamoZUSNXzGLxVQrai1es54cP/Vw7SrNnjEfhWD6sq5VDxre0kpFgWA7
sKa59hF011PSXS/r4Njx7CvPcmpncKsuOHhwxToymca2C5qhnNju0R5XAgCF/IvANsTlIUoXJSxz
m2x5ykdkS+cjztlEXBNrZcMx0EL8Mzbldc1Sfs3lkp3ZYGlpewJ9Rs1Vdp7SBOwza0ABd+n8LQdd
2qHI+lD1XU1KD/VgfeciP4b1kZaMil06QlnbgXhGbjONCqBkPOBK2qLTPpum4245apcchkLHySkw
m5XQRooeR1mSrTUDHAtNIlomNUaGG3l7kbhviyZ9rkNQ/jXo/tUBDhpucewfnD6Dl2I7h+Z0qPGl
RvcLZkujkON8XwO/+xXXnpHV4GcSNuOHmhrXGl4JNXkPnir/GOQj5bCVCKSCe6HWL3fJYmIxKCII
PJQLIQ0H2r1krguj2s4bV+Axu4o+Zvfv6CW9Aa1MQknbAcuPJj94SOSj6ljGAJm4dbuclm9pDqvX
U3q4FMA9J3GStvVVDEtzOu6Cu48MN9jey6Iux+39sNbX3BLDDdpgW8ZLA2HBPVBeFai2xbv3jKy7
kpIXE8W/rsN0VDJ0Rde6xZb9kr61yC1YEFK+iPD1QzYVl9MnyPUUr5ukpwKMfbsExkCjvFzFiki3
ll46nlS0uTaM+ctwpBxzA9KqfBAq+SpImtu6YC8uHk8YFpgKczlDywvB0wqwPgd/irAoC0q/mAd7
NYIIC0TXJ+Zt3ViB27i6UEBAJs2Flv6VDDmRe8av8mQ0rMR54POr7K/BbLFb7mDtvpgtvFNlJhMD
xGnXkG1lazOWgyO0hXRadbJ2EKJ6nTp42rVFihWecUfC4wy0tqLMd0ZG+Ucjg9bg6xNrJaxTEBGo
o3dRxHk5wQiLSf2OhrYnL7a60E9bUCmTxzKaxSptns9WnXBSHw8509OXOazCRwuqPbeB0ZPUiLGy
nkZjxTx4sTS8G8Jy8WbLrJ57rmx2hZWey3KpwaDdfx2GBH2uHTu8Z+5QDkaSFU3CCqM4YhShBAiL
OCzltqY8lHU4b47rKwiCEMqG5C4VSoNagBrlfYPmWLGcHfy4YFF+bbQHgmvOyUG4SfXVKA5zOBxq
hWD0TR5Nx5OtMFTIhaWtAnfNONkKkb0RHZjFhJask0O5T6l6i2D5zzr7q0/zShJmMypIWVGFVpRn
Em5l+kA27BqYu0wizY89VNQ4VnI4dUQvJdi0QipvqhwU8Z6yW8bcKB4P4gduOQHefO+sczQ4Zuar
IXbWrUTOvCtuU+3pe8UqsjJESBewjQSOt37oBCtSJg3BHGRhNkyJXFToIp25yJDxHLt8he8qcprr
YtoQJG/rjavSBSnbYwKMlJPEw5dV2jtEu2gQN+wVUkI4K/NUwmyBq0jzz1LwGtQXQxggbH6u01uK
wWD+Zg0FButn/nhShAvm+3JzfwVPZJi8iVUopWwnj1N+rzFaaeeTdQoP4O95ZSnbVSYOswy8rW77
M68dN3in9n74Mc7S45aLpv229abPcIoyadoni8wfY5HBoj821Dfp/wyNNRHHMziME2BLqyECMd7k
AD6/hQw5iPT/SuPPXAubiyCVXtU7RSRMtCWEsndMbKpx2SS6Or4PNJ4as5qfJOtNZ36NpQ39Aq7l
crcjOY1paEw84jBv8BVHMCCewts046c3DabTZKEhFCV0fAlJyNhnUD+2W2JhNEiy1EvbGxtCe9Wu
fI8cxXg2c/Nh+fVUX4Mlhi5pvMzSFP3olfgHd6TE/Jw4R+PVb+x9N1I+vSRxU+z6VzFzdGg8H36t
P90do7241krTt7W6y7Gq3BOHLcBjkyceNlZAPJBzXanjzOvVldwUrR1EIEpGZFFI4iZNnr3gVnUz
D7LCnpz2LQGRrxngjoMXQug7R6Q96RdBC0s5VKbXlx1505VT2h2fnwLrnJLQ/Q5xaV+YsxDLYbdf
8HszdZl7QxDQ/OXOtK2e5Un121/IZm75IYqqe3AIEuIhqMNdwxJVMDXfmIxS67FEfwRh3Zf5Lmn9
4fIUMpIdGxdxVk0juh2vyz50wEmzoFIXpw38yn2PKrtwolPDx4+4e/5Kfoaet5mFJYEuaT86ORRK
YSi1LxAzpeLdId3Mu5q4i+ltpWXss1S1xRCYOsehVwqkgwcjp6LpZl+wX6BgzefQRDXM+yTwXotD
IxAzjevdpi9T2cQNn0SuC64Da6lysJMBBF6M93DPdUjzm/juO4/Z/gNmE4uPxf+zPBS3rk1pK4H5
hZhIKcvtVCQ7myXKU3NZ2vuyx7CtE7XbiYS32EIQDJstO5EfB8YVNJoiVq4/ZHKIC89suEM0TfHt
V5N93HxDpQAUDJcr2g7YmbQxOU86aU6r1a3XtEB9k56QZHxX6KMPtDJTo6VUNs97Da98d9hwnF1Z
tIHHF9YteRTw2OhLQGABut/1/C281hR9B2NE9A4GeQnzme5VGMgYNL73SOxsuERo0W4YO7BfeqtY
zMrUNYMOdnt+YHT+3XD7EIgDK9AxrpfqnDsGIlXClLjyrQEni30s+vnY4sj4URdxQaPRgEf4PptC
o6/PYJWjbo5hM2PnrMBE/k2ICmWeqQQ641V+7f+rEXvkkyJpyFY02hd7wmAkBegK4HsFE/zVSB6s
yzJ3kEUjEF6tHfgqjR/AJFGjMBkdJ0HKhQKgz9FLm/I28HLd/bbGM9Tv7kiKzW5E6oGbFIZxqAhC
eP6gO+Qm5zABTZ8xarlS5NS7LRV9Eiistk+iX6zjiQkuAZJuBkhwwG9iTD9urUDgu5nplCsfVEbD
z8f0lNZwxOlA5G/oLHhaNKlI23bGd94nq3d4QtP/Xcc3/gxXi+50OXF4h7QFULQlLqd0eeRdHYKv
3oo5CJU2ElZ9nvvTDmwPxC8dgwrprxCNRRuKEFH+EjrApDWh5sR/3X1g+c3p4GYkm0sdIftUNmCU
k9aayVRUwgx4vNAeb6L8/YD2qAgZHoXLTuZILWwO7WRegVt9ueok7coFDDq9RnRzDV0BJKxBFm0i
rE1PFRhT/xyEDMCKHaLZxLn61//qKY2oM4H1FAHIyl9Vj0V9kHGThEFqOQNmaZFPOvobB2E0Qpmm
gjQkKvM7VDSj6AsUsTwm//29xouEuPNb7dLDlv3xWVGX/zyRyNF0wwe7atKxmOyQU3VzQ2v3lUoP
JH6YH/mnUm47xfLQ+k4NfU9cq1sSmeRjxpWOg+FNdzREvJOJtsoEEBz3ZltdLKtHqKL/233eWkBj
aVkEWQ7KZj5v4CkWadDyJPoIK3z7+eziGJi1HvFO+Nj56SoKP3GWjF2biEooZr9MCGD8GX+iOovg
YX+0F2r2y/feynnbSDaxPbSeeerX+Y0pgxIfYtro5/C4MArn2615HQRbIFncbcVVXvPNaZDtYwiX
ziQG6Lsi3XvmHEVnjwxg8VUpoTNqjmh/0WTsIPsRjbqAqqlaZ1OLFYj+4/u+ziPItHZP6/qBrDgk
/n/OV/fiJqZ6U94WAOXBHLpl/eb46Wg4OID4gh6xfuQYXQJDU/iJ+4Gf7dfi5tpRekvatkXer4Sp
R8S5/feSlLQHhojumWtlLext9s5a9j28IMYGyHMoUThNsMs5qPWvPcvt5wiwhV+RNCy+Q6zaT90Z
wwss18ArwWsC/BS14yOEmerKdmbDwx0TPCoX1QwZbtAoF52YoRvlrBcNdi94v29T1n4GzSkHCYYt
r/Z92RbdogQx+kOQ3cBrptoWOmjoCIC1Of6bYiInSsca+nPVb7HfAUwGbZJci53xhlKGQNIKG+gr
H06U1dzsxzSDPI6cVY9noUgiN8eHSw06IlJkHWh2rZa8axA6BbdfSwRwoi04KgDXSZ3NxweqjPZv
xfl9qj51vW8QuD+dKaOb/dB7HhrHJKClC40Pbe5MhpWfDkpKk8wHwYjxnKHXlegbTe4HL5WAdLGu
7nJL2uQuPfR5M6mY16H4BkqhblpPdpR4kMe3mZSmRv51COshycL2gnh7ADquHRm3hitSxOKakbrR
LacA48PFz1PD54p8pBhPVG5AGbJSUIrjPah/xaDGcAds6YmTdT05/lXZbsA+jy9knJ+P4ULJX+Jz
xa6583oe2pckDCRmnuzNO60u8Z7yebrmUcE3QcwGTpYa2L8yU4dXqRJi5sO2MMMS/+R52pMsjGLg
jppgeEJ3pjE8DkRSl1oUb5Ddnpe/oimkTUU8yC1lREQDLOeWHdWiBgadDLlMV58TTWVWNQD9XxwM
TqqWHb+/YsX6LcwTh2G0PWxtxjDpTG627fnlRdS0NLZLWaOuw87V4SxMIC0A0jOj+E3fsVOjUcfm
Fm1fh8w49vtsOhar3CSdLPrGolt3lI0O0yvcmt3JzYHJMTYUAhljVJxB8S0uw73+cchAF6X7AJP8
sWB15l/35VGqUrqzbr/Y3p/Z4hdbCdZP2DOZ4/X3SyuFnYxpipNEE53y25aeciil2g9kK+ANiNoC
R0k3ub//D8Y1a5281zNvXlHwr1Emupxqo7ZIjjybGOfgPhHd9qn2t9iWtIW6X/YibpuiM0/S69gA
jBckvcj+OD4HzNkdIMl5CwUt8w6yzpTOsf1bX7x9tCQa+pfzagqcTpwmfy/Tkbe2ctC0Itoia6VG
7IcxBpFoGoaCwmJB02e1T1bSL/Y+4Klqk5EjejUH4exZn6s4CiPr5utAKDT4Qy7yBSkoyngtxSmc
00NEqJm7m8qgeWR9RowK7aZhfGu52iTWVFi8ksR8El0z4SwWCkcBUUYlV6CiRQkWNUknifqu+VNa
QdWQfnGwLYL09kJ9AbI3Cvo1hDCBSKH9qtPqcQExS5XMZ60bXbTJdptSq9iLMq8FN5lg5g0QKgVQ
EnFc11okpfXJ8fiqmQ4B1qp+TiixJhhWxszDvHmGWjecHk3D9s0vLOK0B4HdIy15WNqobCbp7qbA
NZAN9Be8bvnrq8yZOOECpfiWPzqIVvKDhkvdhZOaiD/hMNMYT0T+Grrvkpdkl98xD6XOIlqF7nke
+h2CWRA3ZClxgvsXa1LcwdPawWY3pVDQi1J8qMbmsXEh+byYkw2VPjonMXwJ4vsLGXo+Eghl5Yl7
k7E08V3d17QersFinSF8s5djnQ5N7nWHPM51dKvVuXuXisdCwG1dHzKB7htWW2+wV1pOtUm42j+/
A28CyCKslb9dtUog0Fl9/TpdazHfIHxVjKpi9N4P0reWWU9stBEaEkQflkHf5IRlEU1+LmZox/uh
6fClbB6B5/flmMHWYCof2KUJ9mfEUlQFU0WE7CHT5HGqY73PA9ypAYzo6qhQ3QflUcA1BNDTQDmJ
7xEs60VIGT1q5oev99ipGGiEBJhR8/5KDLb82pN/S4lfrqPBgha90JtC7PFuUFU74jX/iOlaC2ii
RerL8UL0rttTktlfV8L/Rh5ZYLWcBzYscw8JROfvoRF6SDGoVoVIhrsJ3vkn15Joqkc7lEgiqn36
96whkVNjdi8F1K8gReGqagYPlpxahKV6hLieEx6fcmGp7DACxmvvznLJdK8KU6s+q1zLujzjlB0j
YXO/30ySwHDBCXpqFEyJVPqwPuxpCG86N99Ihv0V1iH63iJ/nM3cd2osOmeNf4iR7HtkmmUMpy7s
Y4Ry8wQL6aga/k+GTWUy4mBd58dj5i90z9uigU1ZI/iwdPrXFP6vFAoly9wgfg7Ty26y6udhGUqw
hpBUl1/BUI73gnhtToweaibU1khr8H1htBKk30hl/KevmFeczevBQFLIbJjvP0S+tBxPi8PVUKZa
PYboV3aCJ4DUTeHrOSXjMQ91yQ7vQADj0ssEJ5tqEYeOqamybJkdXI0aMroMeQXVUT8HeFuhFpT5
VxIdmucSUaCI6Tt65Q1gAGZ5boL4XeJoLyXoqAZj9wL7AdvRTHZf0QDAqX+yUuyRxRMnvhcDcLK6
W5w9WIZKTOHiARBzLZS7XEn8GascI2pCrhOxbf9/65rg8BLf7nFZBZSUeLu2KDngu3E9HZauFWvg
TCMZTKh0K1/2N6iTvEK8o7x2BBR0g984EwjTsTTaKgGsSPjX25ePxPRhnSGSLwg1Di68vGoZHsUS
ANB+KOcI+fBy5c6Vgcrwtx9VcEl/o3vVUya2lzATTxHC94RtI88b/17n2nsIOqBQLpL8ohs12C/C
vYiM6XFpLF/7lo8MisHLLUa74B5ZGGbTX7pT8SpAmEeQi59pf+tllLlLaLDYHuQwx59cviUfYnZM
zcvJ9sE9rVL1wwVaS0a0m5VnlZ+DdHDr0b3UkY3TJaTQZ1/SYCaO8EPMHEYZ5UPtt4Le1cyyiR+O
zTdmjYX4OTNlnk3L3yqsIEIcnA8mNhmWV1lFDUXk9N6jQxfnH9Ze5QzPRS5izkuKuZ5pOYWk6NH3
/9mGy2vAM4ijA+0YUTI5RYhWYI67jnvwRitx0lpSBtgMPySrd8Hwxh6qTChLXkGVbDwciBgDJxrw
lOEv4Ojo639cG2uRmtlhjsI1INSIDGINsykVENruN/waH0Dn8ihvwh89EptfUB8NwqROGk4B4W6k
OoLmBBVoF/fbjuB1gqYz5aBt6JYtJ9tyWM1f+nNZNIXe10xPzH5PGE9v0xVpLAg/ULtZWnLVMMhe
Z4GH548DeUUZUYxReI1TkthEjv3n4tuGx0K8o7oUrcocfZ/EMDYrO3mG8+SIYhY4PNstI3sW7Lr2
IU2ZZv304QHe4p650+pX5YNc3hh9MH+aypCg/prldfpQolS1jn50yey8AgXb0TKlP8U1OyOhquoj
JM6riKfwGCJU6yivCYn2DlzX43IFDk88u4eDxQPAFnuKO3oHygIIJfkmFsd1PYRCFY2ibksrMC9a
AuyW5elMu770MzubM0toPVbOZymZPg1KenTUy0h+jZJIdwt61C2oZRuMFjik65LLLcadSI3CW5V+
FKcFuH9RGnR1YgoS+aegKGhvbOPjQ6WDaMbDkrvhzau48ZtrVhw3Ob9oru2oCjLNavR08OEnD6Ly
9gQsiacOokymMABQbNi+EW+qdoLhEzt8yTMLMTDc0LApamTjoJ6oHocUjm6OdZi64BZoF4tHfFPv
9ZewIH5Y30hXnh2Klj7sF8mXMgqGJj4Fz0/rhV1wjlMvj7B6c5XksJH5/UpU60hz4GSEySvlpSQd
PR5VN4QaU4fjzn/fc6XOKaPGHogLOXYizlDFQUG5ePvxkT2ZDwjrTJTh9kCx7W2WU0mBcqFffFLd
KD0uBNft/JZVH2ahk99NdHilmjkEdIlhe73BfpQbMnLv95J0c7GBDXlI3rqKVWFtSG2g+Bg+Htz8
uZNSzbty9NwP8J/WXxUcsBbmU9J94cphUJpDn/SBWzJtMThn3ASkrc6CUv1HWpAX7qbYMVAQmkHN
3MSxfnrGKfTYlhobw4SszOZBhaVKF4H023/rkdXCgEkt1Mm6EW8K24Oa7ef4uhRBIDfQ2QwWRKVQ
nTNu3UDKaPL9fRqbTFEiEMCE9z02E6rxJk8kDGGNxtmQmL/c2eD51kGYRcGzHaubo1OTZjBRqdI9
rvsfFJ80AqKTAQ1ev1u+p89tHQOsJQ8Y1B15xzSBJGbFpz3MvsPLinxE8pRUfcmCZyR8k8V7FDzM
3nSlQ26GADb7td3GEp/gjpqvuSkY4+ZSj9WfakfuQOJRJB1NQZmtJHpottsjwiTym1mQ5QNfUX5r
j7jIj6tgn7oThst3DtZk+fd4ODM5AR3/YdSeGlxU8FmBdyp1vrSCjynSeuKtwDdWv4uVEnNvQqmo
ceqHWOg6av2+qzOmRHDuGGzNPyDwhzkU+04FRag4iCSpP6PHxPoYRG7/9vsRLWNbvn7wifYPHxEF
KPqnQmzo17PIFQHnNohylYe/KF3xuHRUAiYArZAE3bdo2M0RH9bLHjWU6Rf2gY4EsNXCncplPGcU
VYK4xy+Xdg+W10IEuuEJgcZFhnRJIcZ9Dbc2yXsQb5xg3A+RhfBhiZnuwVCYSNI1G0RZiNEHoQn0
zTjm8yfcqdiphk+anMNTgeJRZqpPS9Y6EH+IhzXqpQhMeUyuF82h6D3lxhptxIwXSQRKlVaQWmrh
kZL+2T1EHadc+XvDaSGIkdhDRLhJFGMmVOXbxz/O9MJR7nUXUD/vlQlay9i84iL4yjflhs3RT5+L
ELg86+3mcooxotO7j5GlZlzLh3fj1TSHyVYsIDBI8O/FODv9bmEUmojIy5cc+w4B/swht9YW0q2g
3BZ9ygisDh6muAL2IXcDoyP4LC7mgzftgqdgX7mjqTAJ5dA8bF0L+pPw2dQURX/rNtNY6V6oqa1L
ThInsJPjGtYz/g7Hk46kuZb/KMroYtu6yTQyIlGFu1FTlF/wX2+C1f3CUidj1tC0ZpRG4XxWDAA1
3q3h2qDnjttsWI9yuIUx7C9MnLMbNOhrnOMNKfYoUV5jx4kQRvKAARPhSyBRA8RbprefPEdrf+z0
E1BxZaZc05KKXbA9Sl5GfhC/rrmfdg115cbYNGxWCpoDRfHGmV6iMF+Kgl//fSCI76AnqB83YJus
AoD6mC9ydsBrLsuILRZgya5OsniqV2gpkzqPK6HNz8MUI8pNau8lLpirJUa3zjUZJWFqmLhAFsqe
QF3la2t43nlsM8XnAQI62ib7/sPGcklyKcafYqIArSHVEZblbzy8ZV7Exk2ed2P9dWyk0ynrXbms
3EVcmJj96hvqUy06cSJHE2t3cYLxeEh5SZpYpGwidNiKJXGLCiZtpjuKqYFaAg54rmYa7akTFPdo
sT5yPBsZSaRk5Uc9s3Ivarrn0ms8YYRBNN7Nwk5LHAhw7w9B/+utiklEWbyo7rj0P0jW0wIbnOGr
EkvKuDijG+mKk26rgN2ZH29Td6TiezIyzPOy/p0MmwKMjLutHZNGKLJVCllvGFtQieYH40kWxfiN
HxBAQVmUpwS8a5X7e6Z1PEIhHSf4uLOkEDTpOsmO4oLqOysZSR0r2uj+QQUchWvPNuZ6TefEQdXh
SaCUfJyOskmRjwhEMpt8L052c4F96Gkd8SOraMvyV4EYkIUnyIKayfoyXtVDT+3CD1Onw/1wFuiW
rl7ArLf5k0vj16E+JsBFeGHANZoHCy4ac/wE7yg7aF0zkOJcPxV+1glQYeN4/k9rqgxZZIrlwIvo
jAr5IUv/ie5aUsGEI1njPx3XwL8dwz94F9Fa6QDCacexeSLksNd/lo9mkA0FcykWcJ+XSdg+105M
o7XCj2GOP7XZBj9A+jBrgZTmZxJP8AFJE3A1w8PSx/Zbq9VqrNy5TDQERqkf9AYDfd25XzYawabe
8zVZTb02Y3Q2e36TxTybtGfHIJDonSSFDriA3B3A6Di2v6C34EwbXV+Dty35IfQXkY9ae5MdHw7Y
GOy3Wbk9ixuGXq95+wNshzgOnPYNNJ8zqKWx4jzJGtF3KZgZZI9Yec02HgShl+F+sjnASdPrn8O4
S6O6DOXDNcRX83DvFNdhyriHkYUKNqf4R/t2C/e5JdS97MFC5GS4JfPTTPpYc0NoXZTYkrsbLCv7
GPCdL3aFo8iIUI//YpABF2nR3naSelgeniWdX5xoGkuXIcG2Our85QP0zYzOc3llj2WpbuesS+gq
G7ddnx8G88XS6A0kJdNsolbFWFN9h1mxd3NleuYjXUUTkWNwt68AZ93Pdw/Ztj9n2PNldgc/YknP
QVAQMNKnpuWNRtTVQwpHf8hEpI8b5B1y1txyhkMfcZEQSjA6M6MX9QrJGRDg331LU8ySRVzVmwUR
X6nT7laq61tL6oz+Srs/i59fe0xpFz5PGaMex4fNCHVgjYkxK8uo9jDRu8NTmSP4lNM6cMAPjG49
8KjnlRmuwtAw312p+HbmcxU6L/yLsZPtFKGg3sbtvbU+lzFpiAk9I1qhLZHPpTc0Ea/EQjJ1KovF
u7gHhDryhyPiBJzgBQgvIuuX0OWjZC9ce/zsBkhjEcEIy4NWFg5gqAc6GnH7KA2J4ydzsUZ0pZjx
veR/rFRb+7iOMtUFSaTUm7haKP76R7hjgsmTeHzJpFmI9yzWH0BUVzZbYpsJdN3yFxDTqvb5pua+
mzyNVBfqDucGxwzNPTCO6uGi6fyrmVdBLnyNxTGWK2zTuyUUFrWmjF8UJhVhZH6OPZLmpr4Hsx05
Gdpbn4C+SILVgWg78P0fAULxF84oEyee8U7ppfAkS2wiqwIC65SBci571FfXTzzl1qlsUlmnyzFR
2caytIeQtN3337F574mHuRuu2kBdrIAG6lv5jgUG4EDfPobeMbYkiIJsNzNvKPGuoDv4DncwMaQk
JZ3tWagnvM5/dtpH78e7kwdnA/J5EtTTKBdQPOUc6I9zwxognwY6BxPLoWT30ueL7FjORa8Bf6o3
UC1sJXhPESj7Rn/kUaFyfAVDq80y5OMlyHsb2xy/bsGIY7qcKb0IgITnlMtQn2JIGArSHm5KsUxq
7B4fZAhmogACQdSjKyBtN2kHN5FWcT95pfL4C5iu/psexlkuPUFU+pLlw1RtVLexTfJKx4Onqjtf
dkyQKy5SWIFpEzSg7zHKnQKLVU65WB5kTIbcW2CkcTGA3wLrv5ppqpeBuuMsthXIUlbqXMxFnhyN
vNXSABLYC3498oZPTJ0kcBRqBVJRzfeh3JZCckLk4FRiS5IQXhyDw7xGpxEBvRKS6j8UZSwORskG
u734bwbWRwWAg/FU1cRBfxVPpqTclWazlWYbv6FBBV46Yvvp+PkRwQljdsMOiKngZoxO5YFxjx3u
ChG8MLW6lkjV2GlI7z8kBAXdRNcF6V1qbrYGX/4p6TXqlSnfzScKl/Gh0YFTnHNglBXF2OjMg9xY
zuOjeEiGuhOf60QcdVdbIjEB3ajLyqQWYBjQnsyxjYrGu5TckMwR0wefYM++AHDUojwwQXN0GbLU
UAdhqhtLX66+zSBslqTBE/Z8HsJrgPObF3oL7mXV9FcTG7SkOFXLE6fw4LElxS8px86cQdWIsyQJ
CvrQZiLGW3NfzSupGHyR5gTjPCmKOQJrWFMkkw8LhE/mJ6P4pYfmj2+HpFAdbzEJ1GCp1THgPNd3
xyNScV9qEN/vbcjWM8o2MSgIgWmkrryGwJjJI1v5G+r4MTvqpVTA+DiC90CPc3jIbMAJ/IPk/ySg
eVqysbU7IQ5z5M6BpdXobGUFdLFaTfVZBSpAY4iV0tBs7pZ1h1O3FtvciZemDs7XihzR28mNalLh
Fj3kst7VjHZZQFeXvJVdqQYbmL21hb/m9NOZy5rHXzMZF7TjQGVzpPgKHKH2FKzao9mXkoiGZW36
IxtzqZRHLmm1ZMO6X6mxzcxFN045ghV0l2jbzHw6oIZV+73REX9hQEtVgFNFZn6BxagCzD/pEsPN
T1OsIEzuKjoRb9DHZh6fm00zpb1rygemT8IerjNucFIBbtu8O9hzrOIgVoS6v462QlVEhn4aXsHa
s852U+atXR99ZW1hTOBM4NO4SbskoOmniSqkRd4yN3IF4S2NH6BQm3UGV9tWMW82TLdM6gA6PKdJ
pl7GBnOSPsrQ0usokMRhe5OCTS6rtLSVMEpp/AyBraUYrjSzDLj5DeUIux6ckQCiADoYjvgFhGDp
zeayL/6jpew2UDWAMrrEcifp4QPvZON2Su9GRt7Gng7dXECZW3sEIAvblbljLqGUxnqO1tka4KEV
5MHPdAvHelgXTwN3yvnVDMrezy4r9waYUw+ANHVxGXvnqahOfZkkWKTj9ayiKytfQeH2c90GOsqM
AbuvK5rg12U3HaQmXo7r3eqOs9nD5jakxQ21yNEKNj3imD76D6zZj6Am7S8M/fq5EH19rs2koDfH
fk0kW/FQ3opgoJcfJaZ+NSI0QhcC4JYtQ+VbYVmzKafvUw9GT/fbwu8A+7xrtdtkfzOA/o06ifMe
MyV/9rSV4g7GzUhrOj+55O9Wd98QCwLx0SOko9d4m2UXgHrBP3vI8fgma2KflYBQW8P6ujx4a3Sz
2TBFA8jshQntJxvTqiOnvUrTGeU0L0so6jTG4uUt9TQKDWeJDQz5qYzP8b9NC8yLjsOPFyZiEvta
uZby5Sg36I29UYPSsNWQWMlY0VG+av20wttQHJsIuqh83VDsP0ybtp/PhSOwAQHc3Bf8UMmLQr+K
fgfAy5rEEsquDo+AuCM4ZdKrrevVK4wOd6iDFL81D+qmYLI7LR//3DFxTUt5AcJYoHtDrLq6UkH5
JuCtJa/IodIjbmYBAeONTUQdUzB36+LHjz5bE0CePAcOSXmhrmN5Ami4vgpB9fwQ8tJOptMT3d6C
5VMYWjcbY9Tx995Z0XpuT2LgMvOoyDylgIyrE3pmZYwVTRIdZZ8YtEHnRmezfAHPl1WL7Wyt3aGh
wMo1nxq2apPXG37hwHqfW7GIm9XK+rm4rWzxuuGsdX5FCpw0DHSOsg/zZc/8Yud1Z7dW2aQsW1vp
ctFz3qiWzIwJqVN4bnpvcgineiM0PttjliwSB+cuWehgDCZDzj1yk5rsWf2nHn+W1Nb8A0bn0OPB
xfX3XokpmP+U4tidiResgGWjJqW/yvU3edcNh+dfJFbOyX5VS5XGbGBWICqi2YNTqejiGsAg2SKH
3ByuTvsEnsfp+bFdgPGliiP8QjQNVPEX1fz1yZbbHjl2KK0hgNjLMo66pouGPQ47L39pBTP/2gEc
LIRHOrbXjos3EnKu0dPVqbEX1Zd6Uv0qc/a2sQLjgmWvCW/AFRDOzMy0u3b1B+fu8gZ1Iy0sQNZZ
tmmKYa5Py8E5cpJrKKoKHJVJpD092RRYco9QZ9kP8Te33ZiRRXtiRUqzz1OpkNpFM0Q7iAcvccep
9pHMR/jY1WX5OFo6QbA4lDs+mF4ufBbBS191IIYnTb/s1MZ8WkikxjZXKLaRpudi1gWFJ/VFeylv
A7wQZFSAbjDNR3R9fZ/GUXKdgttG6RJSKl8dNhLldpcilrLisAA8DFvAMona+9GFrhLezJCibtOZ
2OIKmKZ05SMsHyHDxRCIFnVOWr5J0Ngx1yEHHD7jJj0zr74mEk8Erjraxb9AnX+sIeIiTIGnlPYI
yha7CM2eX9EhAWzIQBM1XuaBSX7Ka0UQdgFmXUYnWepbi30+iTNTtdaFe0xabxO0bGgfCuHQoAXD
otRR0eoKdA5Y8uTXFQccIw4tYNOSyyvFphQybeEus1fGKZekiW+jUX8v3Lum8NKXPNsTmvqmfhaB
80FWyEgGau5WMmmEGdDQ72HooJMtge1AovDtLbT0QIZlEJU2k7Xq7ULRDGrOw/HQcaXiGrMKZv9/
ZfKrHYgh3I0iP202mFOyyMESmnugjjGW+41JiEXVtoewiPljbPNbAmT8tXmvPf3E6IZe+AkPyfIQ
9yVreYrOHqeg/YhOBomP3oO3ZGH0/l6EgkoLG1FpAjRFpMq3HIP1uwVbRoW8XR7VVeMZG8OWxPnb
JKeQRBmpsUU8oHhEkrz3oJ5HKs39Itxwo1Wkzt/IlWdfz/0OU3XNUFTwsyh5tXApmA31qVJyTg2X
5xypP12bXo3S61xFG1jSA0lH6scI+DPpimR0LPgIYSwYcngeLMQ2mUqsOFaO7yeyJlWAp83pALYc
77/OLCKpLto16/f/mDinDBZvknrDvuM7+geTS8YLjLVzFRIM2XSbiwc0e7uOHLyXrPIP4xNNNSWg
SxUlGTZdym1KHfmj+lMzQuHAhHIyOPbdwfulRf4/1hEXcD4pU3I+vhnqu2+acc28XEorM1CQKosS
Dfr0I25gRUXlMYzHQsgo5DXvFckW64kuRN4GP5NDodJU3wC6CK68gxPcyeUEpBuHqDwFGjQxjeGK
Ekwm0DVSV+kmF2Mp0xdFowJgDS4TVqd4C/kcZBCUZimOWFizpr0K43uIwQVDhTUGZed+f1P2Xo65
87Rlp1hTgBn3sd4CmAbghNNdyOIWCLRnO76O60Vsk1zkI3G09XCv9ec7zkx0AXDZXHQ3KwZ3NqI6
dGotUInxgBrPO8EBR+AD1539LdzTiDSD5FG78lQi/FSoxTMLilNLTn+xxya2/Jur2EiRB44w7hrL
zm4CmhfR3FqoYloDR6iDYN1ftuzGaOJdaJM/e84f90rtOOZdAgsm+GmN2VhVD7GOWpuChsFaNdHi
VwgUiIFaq3adJm6YtA1oqK9Z87N3HCIjBy+YCprDlzOwyt9hUhTZb5IzKpX+gvqcwTPkrLwfv1M3
NDNVNGNSXw1bE5Q2fv8cswB7x83gT4eFO90Y3wEtMFQPKb78CO1o1GAr2ENyEkL0irMwQuH4LnFX
0mRG8mdeBPV/yKV/1Apel8TPiUsnWacy34xlK7Tyo4AezNLXvbKHNV65hcFsRg/+PMhLI2uiu8RE
WHG7rCf4HYf8YFA/EgkrxmXf4xYnbsz/ExpwzLl4tO7NquTi2jjJP5TXd6uC16n8H/nSU92zr6zA
CXIa9h5KHk5QWWZlUsgqFsd29bDF3jzJGDjFteS/Es7chNetjVya6e7hfUXfQe68u/4pkGMRCMeU
ihhHcYj4fBoE2Eeccb/UkqrNnbcMW+28d4BEao18JS14qIkqMS83I1oKoZLvYZl10t9m8ozdCFOx
Qb/oSwj8iAoOI4UpXaiibcrHqq3/Rj5/gbEuBTAKKWxnJp8lWaIDmfktemJAlPMpPBmV40O7/zEM
savhaK4nnKV6ytsyF3JjmNHEhdvKjCF05bmZnm1ny524Dv5eJCb6cQZOCbXrPN8e0Nc7wZu/9e9r
qR68qsWPullXUN8DoNxFDS19QFxlFkuxVRnX7o1Lvkt4snrp3LIy/Yxls/dS8TPKAX1Om9uit+tI
e5c0HKktJDuvBwoHY9dBo9fIx6TndCX6TqYqrw67xrPG8xKfRPuz088q9sPhwUdgvUnphyedFM48
KZYTqIhBpZtAgwypC8qg/95yrPPrGz9IX+kptPZd6pfPutPD8oHiHod65iInQ17j02CAYAIc5bQr
XrXdjGPmpHY6Jirx9HDanVAbLwsdGRaEr/5dZfsWTs6Ofh8wGDviOaOtrxhbYgPDOrR5Tt3u/e5O
B2fDkS5mGHV/QaUd0SUiEVFDI8rem+UuJ2RE0UtHtt4XiLM23MXER+fSO0vQ4czfKgYW378+o+Jt
vVmgqiZ8l9bBTel3M4AgwqBwHTJJsYiMq1UqJv/aXDRqWmFRNaIJPJkTmeegoMp1LRT1kHD0viri
/SostOiqHVwi1jB64/aj8Op2YnWV8uPH2fBkcSyOnrnsHcoND7FHsT+Y64UKqqg2JDtiesy3z+wO
L/8Dmli1LfJJteVac4Df2uxi6/l3f8BrsaRRHxEIX3LdCwc7SbLHWb6u5jrJ6Yqu8jVb3QEpZmQj
IZGRLekDboRbz3Wl5MsJL3tgLJaRkZthfoogq0i5kIHIQfS6P73aHF136w6Tmvi7iRW33m0gKDlz
OtnXkAQn6MBw8dG4V4Cc1WrO3hHJ+P5mq0J0tG3aTHag6S53/Nj0U8TqlYp4f4s+/jiClYpxg/pz
9gp/ANsQR4IVTjGAXimHsY9l5szhxDu+z7v1qJeqUGeZCLbggOuZzea+dOnBO4usxss/vWLAQU/C
8H/l/y4DpHTR3QdVB18bqis1wrqEzqpNONOVrK7uPKMREDc37gc0UpvWx/8Na+YvPIhlRUY3RU5C
nd96soy5LNKJu/tOtIJTdEXZblBf9e2a/fKX0vS9afc6DD0KSt0D0gmgHiLmznRhqQ8eBziTLw+P
uOLDrVQmALFMCDmOeUuPcQM+XqwlhGwzGvcqRjf/BMPVztXOvUQjIaasLaJ9JeWMVolXhtkE3Ggv
OSudyOJS3pQEk8OptZ3Od4WwilVBofzPHmGqVE5Tc9XM1DcgKLju1NPfTGeu0BMGgBrxFSSwhQ9D
Mp3V5JIVr4/DkAzgEwk5u1jVkNYLd7JumhJFztXR2v76Oc0nh8OpX3lmsFdEET/FIjHWFWRLvy1d
Syb/G8P82+KTcgcwrtzf0yjUFH8isn/qrqPK5bn8zpbbAJf8oFCZuw2+gQuYjG6p2sf2MuS/9y5u
wKr3a3Z8VFcxCt2hFjBhap2BiK7ShZGeEIYq02Gb/70RqTFcWvHWu+nwOAVdv7GR764HZ8fN8sxY
8A8Y2NteWwBIwEsNsyOwf3M560+OvUi8NKv92ik7thJpBwXaDXzkh56+8ndRpycQBfV5GAOUkCVV
cNxkfEXe20WbmH5nLGkz6lLOlBTWNIltutz2qwoCFs+jRI3HpC0Kp4aiikvYNOwfU3jx5juYl5Ft
/W+BwZfb8HhD79SB9ykSmWL5VxwjTvSWHmn9XAxBNVUCZh3P5aK4cZwywkZwEBlxE1zZzVQoK/YA
a6MKfzoizZCR6GDvc8W8SrVoy0wmx8BLflFGOODhuqQp23Kwf+yhRjLWCtYTxbAcHJtioKsqTRLu
WmVLfnJa1T+L1iosXhw23rFunii/sZFESnmMntI6z4FJwSQ2zFsT2XuVB2gFMy0Vpzp7wobhGKvn
hMD2VcnJ/veSELODSXPcuM6rqopu2ahU8/UAPyMX/AfPkMMil71D7aqtcIJdHLbDtziWwt4Bx0ns
BTnAfjl0KkzKx1wKxnEJVt5r1nuDbxc7nksUvwU+R87NB1qTE3RoYvSZPk+cDAKTaBa5PEnG/uve
rGfKqMxkLZgH9mP9RMHIAKbJZZNyTOC8qaEbwxdRnR6cPpqWF50fQS3vovfVyo7vKgJKXDpMC2wm
o6hkAZztuXjKWZ1+CbT9pjPvRwrsx09FBfzaORcQow/o1IOKtlPsoLqNzhh165Y12AqjE6wBqvEB
Sng85bjrXlJ9KtPYxkoBNyOso5O/GJqW8TzQ/DtdPOLusCZFfLfgAwyMlcyADEIfpbOM6UNzWWUg
JjgaweI6wN4Q+IuK82sac5exFO0olvO6z0rxHtX6/DA4ix7Goz56UUGNIfLbT4wv17QeC5kWhQcv
/ISSuUTs67vBiKM1rl6zteyYBqyt2K9uWXbt3U9DONbB2M/LvJMPmMZepiU7uGjv8JabyTKtxGFd
qnJBmT6Ki0Yc2ovrX65UQy8arVl1+pSIFCNWVkmkxtNYMS/IWFPuqamQ+5vIoQsIPiuPCAAy6X+X
G7lhs6RYIYuqUcUgr2HqaaVYmqExpMzIyBenRqzgr2ARELU2CcgS1BO6erjpFiuzNp8YasEcr63Q
+eiQG3QRhfNTEfB65y3LWIFOPTf9Lu0mf8MUrC2cDSdRdWNqFcjmj4p6+iAYY8vD6vtMwX5uX6DM
bL+7BIuPDA2AflOTVp5NfZO75ys0Cdfr/nKzHGeMXdFiRMF8NbSeOViNtPmFXhZPurnlBY6jBbfg
c7vTwj2a2Q1nYFKHsve6aW8RYPwpjSjB2kXtR016RAqZ2zF0Haj8z0m1ZcbJaZEyXDpvYTQbxZmZ
D7VraOLjP48duXpJLOULQnkfXcg9K5anZ/4WYu65ZeP1dZNiUa4WBWwZ5SZnggiBjMCy3SOaHJNc
tDOqMYWiuXZ7zUMK9eR51ej9k2mgNa/AvApy0Czq44zLGgOrxMQNH+YxJUyfMhCmWbwgw/UEbFgm
uig1L72+oFGssOJT07YHH2AF9q+xqVZEN0mWYvqKYLpj0EEaGF0JIdDUbl4PY5i4iru75Dj0rT5O
6mLQdyH7+KVCeZInUmNo6YBGqVXXJcDGlkQOhm4SZDNQY2fqQuHx/DMuy1Wll9HslmoCanYzXM2w
0eTXBCTbUely/286NOP4uWxFGELDqlMPdVbwDoplyPPW60oPXH8GEsM1Xqt8UZq0nzdVhJkeLQjs
q7eaHdmFQOB8a1kLC8lp3Pfwf832n4TYSE1oWLDnjW3LWxRcGt5Tk7eJ9f+7K0z/YrIkxTkhMpaG
5DUhHPxAGtVrL+DOxmm4zLiXMYLB8KYpe1FBE9b6zmoPyRi/A3e5+MCJTh24gLn6MUmHF88YQrTS
mWlYoPxE5D5ADpx6dLXHUvYtnL7UAUJS4f6PeCuNP/z+F7ul2m6wPqbtUIzAEKxN4BZAilZiXSop
Z/dPPCuN6GokIuGev1btitVY8aqF0F23rSYgbYVog2crGF+3AdxWWdyZ9BWpQlyQ4xc22uswp3wC
t8MRqqw2MAo3S43vEQygykWl/sx4yH+Wdzbfb5ImTXbmqQpq5cJOGkqtnGtQjlNOGLb+b+k9uXKB
CeT801uVMhVHkZnjIPzFiv97en2Pbw4dWr718OrLnfWMQUrweLXGa7fM9TY4RDzqENEcHhAElqj4
Ssajvi5VippWmuLP1Ryez0xLEft2qNI6Z8zUG+A8wH77FdQIRxJsrXRc39ejy88LuapsLZqT0ebf
VMIBeY+YbQEf2oWiJzmkvKTOeOQFmDHfpL+3ipaJ3q8I65PaDZqphzDDyOlhph6Wj6GM+SJ+CJnh
OoSxw5cVhcdAZErpwDyhQWAU0Fb6F3TYPQv/v5S1kBMDXwGj8zqmHwnQAudPHbmxZPZqCW8CzaTW
ROoeM4c1BMZweIYr+s+H8PJeg9z4gHe9aA3FqbeGEL4G44p8zHL6Yu32Yfpv4VoNYU9Jvl5rvvMa
JsvBhyRfF20RHz3Rxa8KTH7V8Oq02pYpGkDJmkqazviX7FUB02GNWOJ8aIIQr+VqPjVAejYOk2R1
iElCNIGpRAitAuTJ65sDulMY7dQkEdJ4cy7BRAnArSxpnBGx5EQllVT+QiacWKy6faitrZfhXgJl
itSaNQLw88R+Rt50zbmK+w6grBRdcFvn6vAJO5oyMYZKJvouLtc2UZKPlW/8row3OYnBgXsW/Mj7
whnwXgrykwyhSUa2KnWBCTcJ0/1VmGlAH2ABJZ5a0mqaRuipD7UbyvR16mfbWXbryNRhDzyfNm7p
W0SOxC3qOkS7hSDsYCDAKgjLtALM1DmKcHw43DB7T+UlTBY2AZ2BgtMpsAGE5rLv4kbgXt22HaoX
G03Ah2MplXovqyI1bNLx6UeZRrNN3A1JHjiGdCIB84lOvIaUDJLE2GkX4p2q4I14Jk9/Tw5QjLgP
9NvCaSD++pc+CWh7bnRM0bvryY/X+x2DmZuu7opfptZPKs4a+sHu0ZUrOoWzFDxorL5Aa567Zion
rimonid4XF6+UShllvHbSto8sK5Ymrq14qYKUF/ATwBgsbzalHbKfoXBc0u1pLLKDQX+leA7D0m0
bLtIcwVmQGKATTUSkAIPYO5MUIi5r5kR4ZBjOMyop4Jz8TFp6BCeQbeB8qfvG3wsh1v6l2sj/rj4
haikwZw47Q9sUktOBScFqgdsKapG2e6PXtLybAB4wYI2pAbZChMPfEEOiEajoOvqZ76uO3qke/Jb
+7TdlwGML4ClZd5sJfJtOiX4noD7aYBwNCvFVBKP+wSPhJUrMC4ImNqP1SKDKpNrnJ4psRADMLSp
mh8UC4E9IJoUktMQ33Irl1kzl8UQV/IUCJU2yGuA0wKfaGLLhlBph57GffCDxPNMiDqJThQKSDi+
2+qGhpwP0/cL12RoS8FpZaJpKMqMQ7KOUtAXYIHFexFbv6TgS6S028ASguo0V0q2NEOXxDCeTdsu
EaQIshGfU83rnWSzGr7VrYoRKUkFN+slmZ1KrOqMClLHKn78wnomUvyeAKMlWFtcNcc0LWHXiFi/
N/XTcV4DXJv58qIvbWSmHZ3P1ANmMQaD/AVdFkAaYJErA/zEYQrL7XCsXs3TiOpoaQIBDXWGA/y3
Rf2PjQic9G+wGVSUHpuWKa19l5dRXevYmR4BvSEQZmdXjV+xaocDZAiL3w9yZPevNGUI+zn6SGDr
xdiu95o5jrJvaA6tX1CCjP//+zytFbX6tazjEEa5EVDal7L4UAy6gO/ToByw/x6dNgfAzYdzaLm/
1HA0veKHM8gD6ZEmM6gQf3cB6pCgPNFBUBHpTQ0i8DOafwfbPm0zhGbKrRLyQlOoO+KjmHBb5m9w
zBvNb32U7VBj45mplwFDh3baU2n+UJ+KMFXYS9JuKAjNMR/YJr+hf0a8pjTjdZ3sNBFCdIywj3EE
Oqi/P03wAvkPuCtE8vrvYLup7S3LWAcyoVwKiHPlSJxsE+zKqlbvx3bH0ma56puFMyAuXfY1/Mjn
Wvpv/cHPTKzW2MipVG6nJz5oS74OM0c4aLG3qm5d11hDgukp31faz63bL7ssc5/s63BmCsCfXVPo
l1P3jy9Pl4qbfxhRp5ooM4lvF4fwZQBQFIcpDBmk1JbrIf9wCXkRBdG4IYkq0dOiEzRdVDtyJX9f
TKQ9lN/cI7CbUvswT6jwpnkPVa3K9urpAxI4IoJ0SfhxgXZSV22/nJdbzRvUdZnrZ5et+VEz5o0D
lPZueTYK1ISKkjvVRST0KYbwdCqjFGYiCftjj8CYFXWc7mGoJEHfegZFF/h1i1x99YnXGZaozyyB
TdVGSCOtliGkIIGd6gea3mXhxr71/N+mTroidm7qzS6Bj0Zbpu206ph28L4JdbgZ45GLo8Kasaxf
dMDkX0XdijJ8B0uPzHMDHy/UKtaUqfRfJ+O63MDnK9VTUQYtA+nPvTx8ZjLfJUvE3RM+9xZbDXU+
0MfqU6HlJtkD3yS7PAhBi41pE50r5Lp0tItR9nYK5bNfQ12ML7f9vewLQNYj/n6gN33j7Rh3wV/c
sIR5Bu6EVwNTNUSpgIf8FSrnOvkbnnF/ajw33TEfKhkfz79plFMAB8o7oF+t1s5F8gI2OCucsrC4
1ikWHcEiA4INr/B9MJxijYJy8neleNLwMPCTKgorfjYGy6pLX3MkZoYykJxOYPO/YhqXHsa9qxa+
sSRnuKVLO+hpsup5lasNFryQZHtIKEkKwm0YxqkffR0l8GNOSuL2prVye/+xyzkvhfG+EOtxxnrU
fIvwkAadFEzP1r8u6k3O6U0iruD/5s7GNvLbeuJ4yIRGxUxj9XmG/ZNoh4Qr4ybPv/pLO8I3UGA4
C5D4mYoTEFVXqa5UH1D7XwvjXDb0C86QuBhkIAPUZ7KoCOnCNKPgpCDQ7eEd+ruWMxaDBZx+bPje
maTCP70jGTCwrczWLjyffLnM43fA8rIXYxI0u18Ri3idS6RGYOze1OdfrCNy0mRe9vPSRCqsnuLl
UksrLLAST1cHGgaieeZVOk2nC9sEE6koieMMuZtpvUULa7IAV59SLZQvN6OEUBmhrLqw0wDoncKj
HGOXsMdqNuEKM9MP7CA9dkJ1L+KRyZmonxLs3DZeilFGUMUAYe55wk6mmLje2ZP5gK061b1p3+5g
y+ckwyVOOJ9LrdRs3saBSJ0vPLvPJG8SGTqM1L9pN0usHzPY0AkGsDXFC4K0ou70mGnt28cVmFTl
1rE+EjZJarPFGCtj2mV5URRN2IZPSiM9hxbOrr82PvYSMnDmZLmYBG8KFqaT+ySDarS01K1/pSwr
7wbxmE8s8Gga5oQ3YGqGZvE39IP+IMf/SzTVeTnKNO9Lo2RGjbZNedPC6pVrRbiVsH79q9saebsf
A2fX8Li9bAV++G6svkwc41dMgbtC9A41npivhGj/FyCDxhpySpIniGNgXApNKbzGRThsVwQQEETc
QLqXI6j+3nU4XXS+NfabiHan2QFINDGN87UUfhj/OyS/t7vLQYOC2U7UE6VYHHPFVSnj8o26lXwN
eo/4y28MkH1z5TofSlCokSLsaSQi/fXEdZHNtf6vxbKceP4wKZJ0hNT46/mVlhumK7JHoOGDaCW6
b0b5lzA8xZlgexv9RzsEJHlbC1wOtH8bulqCnMC1FEU+U95jJ1PyzdD93jDi30IcdkAxXStlzsMw
ft0M5xkehrQAHmXD5W+KRrrr2HfKKnxUZTkFzwntUBLHHRgf0XG+f8vfacRkQg34aWiTna0QoD56
XbwWMUAnJ6zzhIxrLcyWjc+mfu00LArXG6UWT9d4xUQ89+KoM8Vcd/nJ56ZO4VYQ5AMJ16R1Ubg2
gg3/0sn4QtozMTF7jhN4UpRRZ/tou7FKsEXZ9o+rJFwaiSaGAke0usf+WzIvefziR3Ann+wVwlqO
4EMnzptwYitxwZZmq7AT+Cs4TE8rFsAC/z2d6wOXKZGrdZzZRHAJJP1GDYmtg7T4si/0voip7F63
olQfT+Q3u6fl0TPUzZVH0DOrbHzZ9TCpUc0FD2YukHvZisOO8zayd0eTxxccXcTkfcJAnFpUie/9
EABmdrFpmelQ4PfHJO6V4Mpw7BI7H37JaQjeXEMBcoaqAy2k3DukLIl1LDj/gBdGfS/8XR9Ds+hq
mwFlCyDvd3ocnuCJZgKR8v8UhGBOJ+uhh2iArtL7q/h12+BGLGko+OewLBnuyrquCZDgWqLjhhVs
xoGIVU97JKddDPJcQ0QXJXMbRmXJMOnkEs7s0n8KbjL3VSn3nbNVzv60XPiIkwKTS+XHlEG20ur5
rk+LkWinxw0/GL/kcotaboljQ7Z7A35ov8+CDfpVi0u1e690QXZC5QZtRUBGirBwOEAxPU2UyP+C
itHJsT+q8C8Ro39oWnLYjrkR5lEsKwdGrK7mRlS8pmuM523DT2wDXw5GRhaWd+1TcdB3j5EQTV6j
UCTFlPRKVoSMTxqhVoVXTFjUQYxDCEQDlq4Z7zyru6r2AqHcqyMMyROnihyYcluAWROA0TdswoG3
eWLywq2QjHCltz5lYKLgI54Je/0+gha/yTaji06V1E4mZKoFn9DbRL3Z8Xz96FTKRRKTVLeemphS
lLVwrEVmFVDBlB8COe7kGuG14ldjOXHipFV8soPhLCZfvH2kZ72HnV34u1fdobKXpW7HWMmSLu0K
np2CREbfGrlUxJBYXwp/8ojIzQNY6Xsw3zOnXy94rWlkGUf9wqzC2dAi9GCCia698T9tfm689wEK
lHx9DktRc1/C+iqf6Aalm2z7/tcl8gDH95kT/hcidKkZHUHR+2SOYY36oyV32LSs1Ere5zhcHSyv
m2jCW1NWgDeNYtH+bP+8erADZVLVfTwyxbKX0SXM2p1aOUEqEBIRHxaGL+epQXZc0woscJEFGcvt
vSJiW6mBVo9gpqOdzcZQBfil0khUSwkflAtN8Xbv3fzT5tC+pHKbfvwpc/97L15F5jSA55NfzV6E
VKnAkzFR3eUtbsvGSwmdhTrSiVrhZ00dc8BErbetvCsS09GUJo9G9eaD1Cjycygbt9/zQKUePpBm
ZjsyKIHpWJl8A7CGOTDpsvTIfn8ol9LklUOlmNEiHvNyxyPzdrCV/CAaUSO60wHpSPI8sGIIf0Ks
EG6EHA0uei2pkDcaIFb4ZeXMErmiDeu0aYCKf0ycwA3ysqkHNn/Nh6V36hLR/lREOOmtjRHBA/6H
Z+7XUJdsLitF3JGexJSJkjelTCTgu5cTLHCvcOuh7Z5X1iUSjYf05HGH85ZYUnwq7mZbizbLznb8
ZSBB4axqlzyxCk8X2ebWx8XmcTwRwsdYRee36DJs0yt/gpaQochdSHIfMbr9CFz7F2rga3dJV+EF
8d1dTu4qT0WD8K4mF+Va6ENBA+m5EKrTGpMCf++ZaCmvPoyQps2+JitETa5N3LLXtCcwc97qVEsZ
2OlAdq7YYVB5/bgdL013/I0st4Ai2xV1aK2oQzQJ8CcFzH/ejKnknNYGbu+/YVj8BBJ2pPI5ano/
FOJ/73as3SoDAWKfIZU0dMKLa3d3dN/2HsunCrEHhKOT43y7s5ldqmj2i2K9sht0IgwFx5pA8YiS
hM2XQAPF+TVf3Ofibx5hIRNy2En/8jn/XYolAWtfrQqR+zReti+8T2Jd9cjD7fgQIRYNSFMdkd+b
RW2Cy7BbI93QIbQvCcoccFiAcbMCyCqiviQOFOYL7uGOhAWYWPJSSJk6bcUAjsXx5nj/k/viMbja
iBLROtvyti3QnxN4enYpiStwDFdy94TKj0iCUlFlaLcsxD4x23FNqCM+eURFjHrrKw+OI0CvC8qR
t1mUELSNY4FhzLUT1vlGlnqV6KwiVSWpxhj1TWNif/Uooh/4RLPJkyzRwttM6/1zNSOKHhwIPkP2
+k8BlV0UdwK4jo9qzPok2aCpoxYEqRHCj81J5fqIXIjpkY/q75zYaWR0h5lD4GfnJBpchls4Nd6U
ar5D7h20hTjJ3M2ob2sfBAzhXKzJsOBbNHhpY3kunDsb9TWqbo+rbnRJJmlsSKErVLOBDRqGQ0Ef
TW3rP0zuHMA1Sim8hw84PSQs50KJXDY6aEI4QIpU/GCmNVbx7tIwjPnAz5SE+kpUnABQtBQxD10N
wkkQUWmjP0RgxY5aWwsY5EjDGk30B/OW/pzbITICalp9cPAJ4v2OApbDT2bZ5dpa9QKqn460VEXV
rX7ajDs/Bkd1/cg4yA7Dlm4Inq0jy3tJBmnKbRyxWgG49aFopENylc78EykJFqnsQOeDLoXPSSPu
NJQNOkNWMKzpVEomthVYtj5f456RBuhyRySzHaVGxozhnhXRg0+V69kjCTLQKHX3hohS+QDST41T
hOSBh6dy6pQiYraVJo4cYx0AQ6SMQUv/WvcAbsjnQVpr+iW3q2qOEhNdDk0QlWCcSEMsKkVC7TXY
WDZlx/pzJcI8Ap4rT1tCKNrTeT2KE8fviX/XQqo8y3EUWUk4m/5o10esU3MdH+Ckfhw23RBQQEJe
UHgH9UMu7f/gIHChshiZ8M3NYcYs123jZwLPl7hc6o1a74u8MDkkFL/yI/2yxcWNiUw2YZsNoNAS
nEZ7jKnQXHjoBiWB3e6/2e57orqTEfBpEWc012OR5esb5fVjcwegI+bpIBxLYQX4P4gLp4Dv5aUr
B6xVJaiUbXIpJjCzNCpK1TUTdY3fMqeHhD3VBAfTqOF8uBXVmlVc/xl+jr1uy1qTXCk+BgRCJQt7
qRd+KPA4kCclNPes8DauT1rFHZCLV5BNgIEIsQkIFquKC6EffvnyfrQVVtkqEbQoFh5OX20ZXuYG
lXmhT51PilyUBxh5THlUvlT4xU5BU8hWRYMjDWOyCstDHPyiw/Vunwf7n3mTDJbZrh2/5RqrNFL2
uwdDGNsiwjJ7WEB7U4R86H7KWPqHQFbXbh0g0RIga2ata3dO5tyi+5bZEdMPaazzXfb3GJdajp9W
VXa3HYKB5DmOXzpArcajRu49hidiJqJmEmzGcLnbQaM4cTGoUbFdqwhqKVjhEJv2lLKrFFNnD51m
Em1h/Ne7zPmQ2yXDHjKhdn0MAdVeO8JrqevKQy7m9yQ3xMbE8fu4NOdn05Sg5dzhKb/bJXmlSYaN
ReYMf6oZb1vnjdIh/cVWsuGuDuJLojIAgSwej+YKCIaXUrfq2nO/e/G4kEnf20diuYrCd2XeuOFe
W0ow2IOtx9Sk//8vHUr7ndUC2q+SlrMVFj0uHRqtWNRP4Jz1+dV+utgKSxOHR8Y/QJ1GTzqv7K61
5JSWUS6sE6q5e6wnfPztxzunYKmvRk+owh0D5l1xxw50RiM8WPipbWvEYLGwUI5kLX7JtYAaIFlm
bUfSWExr4Y6wHd2iwqG2e9jJK3s2A+u1WLWNp3alTH36//KIcIvvIBQATtl8Tr8BNK2T0ZlW+op1
h+HSAavm0Tk9numJaDUEKwrohf++RohZPDQSBsGBxsVWOscgcfwOAuZcJ+wO38FniucQMLS9mQxt
D8KipN33pd5l9WLoQsaYe+4MlAyGixND62grZB65rH4RCnfY+h0hQ9Dx+I3ifda/7QFj8rCyrc0P
KA/sJXxlo8fI0RqR7uGB3qnS2ukteF4cJPgeqPKU+xiuQr6jfAHwFfiX5jsCwk3dVMYBPdD6h35P
ts7lVyeKz/pzaHMtlWlaOdBZwI1oMteYZEhXSpdUTHvb/14pjoZ6YjkDl9vRKpYIWmCf1Z4/HVFG
8y54s/Shw1HHoRXe9cXHZCuXgEjnX7/TKlct1NKROnlDWAxsNptbDeTo+zR0uhS8pB8vJzIlt03Y
pMKljMtmadHia5WijxRoICdBzAM4PgHMyGM59tdgwO1cbRUCLeK6eIquaYnUzmjj3RP/3IudT1Dg
59hEU9UU9a/VUIGKXWpoEdAqaCP7nW9mK2eJQ5BoUG5GDOi20bFhDzxIyD4bJ05F2jV9HnuW6G4r
fRHLuS3tLmQJX/9g4XuJqS2cucOiTKSp0AqrO0oJ3Hf0XdzVrcGOMPwLPK17YZIjyseYAoaDkFz0
D8ZsNgTvjnB3usflsYgC15l73mKlqJZ48agjoynh+eb1W5X5+7qWxQ7CJPDpQ+NHckCSCSuzVl8G
kSN4uM4mDGHdabi4Nfwz3F6l1vTCySkyNdvhBX9itU6TZG3G5IvfCy2QgDhMwsU7zG96zqxGR35B
Arj3Oh1+FSv46zWDltP3hPc9Eb0c1TZ3X7oQeHB5AwYRzYdTW9I7to9EG40VlBEE+oKGe8xIMpqx
ngTZCkF2uzhSVh3A6/l/1cncuxAM+cN8/B+PUa9Yp2ZXgULx9qasdq8G6pejvftomagY9PwwjivV
4CKDKvXN0BcbRUH9RwteFfDlGUdux0Ak7jvVOA6X4RYXD5GHebUh6PtJ/IqPUGEl8Gxax9br+DG8
sii0ok76Z7O6RXIojQLLkj3UB3ulZy9ns368Rubvblx0a+7Hi1dw3BEVq4FjbIZGy1ejnZAhP+O+
Vwv1l4RBCNv8Cw286uJ4tc5ZigKtg1Wcv5duIYv5hw9+VvXP4gPGPtBZdwvD8Zyxx/aOu+7OnpLP
BZq1skbQmueUcpYUmXMfPNYHWcsNzauKGg/ff3A1wgJGvPsHw7rIyBzvJlCyd/7g8BgcUYXu0yvk
GtJsdBsOn3U/vHBHYbPZ70nx+Fl+2enreks+Q57Veqs66LTsWao+X+F3dgyeNABk1It/JB0vmKlh
cKH/1GB7SZT4ypRB6ssvt5tFGliP/mTwdMHxPi/uDDV6NyI2diD1vxcVpndvpd0/KL7jkLUmg0Q8
s/4aQNLcBs2z4vdI2W3ChLWHaJJ9IcG3+tDXsr6a+zxL7vPLdrnaI8TGYlsR6qjQC1EGraUnMkFp
vPyiXMs07UfFscumUDsKNwdYU6b58A1yfSMYlUcZ2is/fyC+6i0puAMOuDxnG07k2cFlL6mix7qa
Pn0NhPy2I7LmlXu/VgYQwc+zeB29yxXPpeHTHjBBhwtC6aSx+2mTmlxMk4i7wgXWNVfH2W8GCvIj
ZAWKDfjBqxpcscgjdUSrE//FAnGyyZj5F73tWR1UhswfMkQVJn4Pbxs+D9RG/xf1hrHx2se+RAvO
bdzriZKFr6xHw5cS9BneNDT7z/nh/VQnu/YSF9GWPUfiRFLoN3yuh8yxCKLZIHcpfRqrGHqVwqpI
Mi/1FnGpQqVRVbH4sIxTVnn85RnBOqeknCXS0iYJeYrIRf7SBJCxQo7jCwq0C9oMKZbhUW8ANPU9
gyd1Pv/Bn1m1ifSPU6MOeJu8sBxmvtVgvJ25OK4iJMRdYD1ufHtSFYykFvL5Y4r3RWi+yjOHaTjQ
AoU7A/VoNIyjELys1LH+j1jIiy2QtFvPv+DbslRjDrYARHrJ3eCDgEqF8ljw4So9231r1QbAWmHa
N8XYCCqu4bWD9TqWaIJwR7Dj0KSiiESrVVBA2W1E4M5oygPmM3c/PJgXe5txYc0DkNGoWB05eylb
YvapMn89sgx9u57bXRLaYE8iWHJ50DZhf4BYH8LeA3NOg74EAdy98jpFF+hsDEEvT+VAt4c9HZFU
P9rkIL3rFTGx8r4rD0mX3mXKlrStav5kiV3ko4khMmxtTp7mDjhpCQO6R0LLyb3keUPp3njJ3WBk
9dm81dfeXVvnl4bC4TkaE9xet0fj9CuXbk1twF3L8flKbwjGATcpfmJQa/NUh7tFBzooEx7bjHbo
f1kOYkjHRjGm7J8QCmGlrRfOx/FIf3puU8BgOmtzulKfcVWbpRShyhOESr/lB3/Iu6bU82bSlMhk
NSy9w3x034/K7dKM6hjuHe38diKcuEWfCGC3LwDeL2KETOLKJrm3ZmyClB3k8CHYNPWlNhIiCP/B
B1vmPAZKeQqHBZfLC2CNcAG1PrcboBfVB95YTWCxTiPHUZGNmFODEu8Lyju/2nNhC+OUNlTYL6Fn
8U2AMedlInUgea0WUkqUwqmQCv2ClwLYL74JvLM5hZWvlmmn9ztgMi0L1S0HEw1fvaPyZOkmOCoR
jhQIb08ScTGVSziFiJN43vRf0mTRsBfRpDXRXA6JI7alVKkfl9X/genmIk74bnBzs4/jpjCOjgl5
dMkk5+JWGOUS9zMo/SDObL4TCcXigcUtjwOn/fmYWwdBkyaIP/Hk9bmRIPPVcm4w/5nDM8dCSUbx
w+LvpgYSpmqYNiiYB9x/ROD/asDW0FD8Yl+Zf5hEUAXCbieLbeL/FaZQ5XLGnFNyRml5JtQ1H2cK
rLTJJE2RGALw21dpDANrDuGnqOIIlKiP5ePXnzXkylqDUON34BbflviFVy9EF0AZ9aQEoOGhE4/S
qzWw1C7PLhrJ3XxTQri5CBuK4LlV6oL5fftPalXW5SQokCB0iG+8IQOM0xG8bho/CtGzZdyfKl3w
ImsHUevzm8s3n6ir4B96VqRSusS8uz8rWORK1IC6FKHuY4ZjzZSkpY4YlOebp20hz+Ctm9PjMSQ7
d777Z+fFDqgJdjPNmxkJAepd9bC0SPptbIcBwbJ1eykbYKudjwWCfjfrNF9MGNNoRIE546iSlSWC
CcPWPQOZlERAJKrr/fb7tzFbzXn5MDyfK8ZCxNIBKBVkCcdH564SkLLQgLaGLoaEmH1TRSh3qkcx
27x7D8/actmX3BtN8CI5KN8fAax/XJK+lwpS8c254hRKZhg8qD2IupqoRYy8IpvvgXDP4isTEygb
BOiVkIc9quwcdNQ2bxXPOY6YHdQy537gNPHuAjayXU3am6KpJk6iHgJv4/Uxfc8Ju0Sk0JHWv2kz
DeT+RWiZzy6F1q20RAX354AUxkW1rXBeMaXsN4egAizLiTzPvXgxdeZ+Fq4qaQQX/G69BGv2jISp
Fy4VWow5Uj9FjMaoGa7rKwMPXg/oy81uJUdxYWVQpX1bZ7sTTbGaLCCQcrE9dJcDNfYIxyyJis51
WVCT1UcVPgN46qSHU8ESTu49kh4Fk07McuKSu0kOE25obHRL5VlCEwMXK31rGOiQrKmKkCMb+wqP
Rhuy7J8CH21LBKsi8TU/5LLhZrCpwGHAYtfJSdZoOgwz/Cozd95J/yWGnmm3Y+Bvg9ejazEfMRTa
KMTKUr9jbZqi9oZJBEc8OP4qtpYq/u9+d9jy64es55RXhk1ISbC5RCmaR6dTMYicob65zdvY2z7g
nCksn08oSQessmce7SENfYbXhmBjpOIV6fYdlCmJcVCmb4SLf6s5nT2whdglqHBzeWdBqin7PyVR
4J6xpw1FAfOqHv7F3ILdOdbTIhT+cNoRSYys0Tx3eLgvXkicbfeeqi892jkiVOjNNeHJZspZKt1H
R8e3FN8emRXXAIs9I6uwM5AP9Z/RRcOswF7+qo7rah6j2z/GkonIfCgTUsZj9rYCHBZ9gEm+5Z88
6PSw4rjLjle9qMp8jBdNMxqBO4LT/bYRc6ZFw+qe8CT7FX8Pe3qotS/oQ47Tjho9BlfLN3iW42ao
5EaVe5PzcSlDp/8T9nLmZI1/G69SPi9bgDUUrbthTlI2fPyn+RfypEnHa/alM2ndieEPD251RoPx
e5qg1IMWV78IBTWlmr8vqkwPypAW4vvlQLH+xyL3rlBQMlO2n3N7MIUDkm30jjB6cnz2ZEPzicmb
wyDgO/SZUX36TQF9zphzOw0qZi7Ur6dfI+sSGUPr2WN+9eYNLOPtK0qMcMKk/KeRn+xownZ8Cklq
h9UsbuIz7T2VWd0Jp8Oeg/0R5jRImt95EG0L9Ln28VYysiaKNTXXd3AlpmjJCqe+PAepa5l7sted
+YITKYSDp1sLN0/xV3qlr2sPxZ+Py+6PjPz4m3S1aRxQwQ+9wfgG9hrjfY2n/jG6eIKyiqPdfQ+/
AxcpxM2SE+bs5piyjKM79Ym8RoiHS3RRQyeL7iVfd43tywUHxDLaNhZ14KrUp00d7tHfLF/YhsU3
hDZyVlgbd0b+x4+CYDtJp2Dv+qz0XZHOAxG//ZW7yTK7+YIFPINyFuSloPV5R3XS9/myPoAw1aeR
/cUEPfqNiZVZl2F6Mia52dcB7cTRgEDmwTdskl3a7HIzy1nX4koFMAM29XR8PWysc9/7c8/6QVCS
UZwxQRixUc4ayhJnATj4ylP/PpiyjSm/qyXhhD+USahwJGdtpVn7dMy4ZO+FhaUUXD/sw4dd6L8k
4GfKA52Cf9WGTAbmntpMor7LzzCLiI5A/zfRRW921a+0LWFO74FawXrhRr06Rf4SoUxx/TQasZvD
gemQGDk3brV0fMLXh4VI9uKhGUbfbBhcCpQhEHhcZ455GDVRzXjTPHvQmRBZRyANY8CKP2xZxskp
kyqVcqvf0fWsAEiZcs9ay2nI5snM3foizhCgxUarP0Gzj7KquQxUb5bH7q5LHMVnB2DyerdtO9MV
aej7rTtuWfC8K3a7rhmbuJMhWxUEORsTuzL16OvfWTV82xRi55MzTVmDkpOLK8u/KQpaiqe2opzf
dyhjb/rbFxvkySrVRyDP1HtdD1QM6+pogdvqLYOTfW5zvLFy3FFPwZRAXWi8HCNhLa4R9cA/CnWm
CoTZMCkKZYdK0aF776vUBfUEjf8tLxYnqK6pC5mEZ6TqhjSF27fxVXcDqDuY6CcyIt1C1sUoAEGn
YJrRDBNiXK2cBz+YuKTF/JRiLyz3kuUUG9+qqLHNie+A8O7SRbBRtHNyq75PDV/z5HYrgBdSSTUm
f3C9wg3wdtIMY+Gj1WPI1SNRayYf4rDksIWAgN2L9sxhqIqAL6s7FxYLH1iSEZUFZ347fckAMlkX
GDMzkaY+4jJazvsut/gdpQ+VY0jjfKyY7xd+H6Swwa8U06kzMQciOeYGONlpjFS1Tp2vKLRZ4fLn
fUoYXuGbDd2bG3FIPdPqUm9QmNr4YklQyY/TiteFBsZC2uI2R3zHGbEESQOTTwoXOcIJ8uqgyq/9
EJ6WMbSLNSOf+pBME5a8B0WUV14FSqhgtkS1thncDnPQz/WzLuu4woVCvlYEKded8Bz4iKFz5y8X
LHsSKX/AKH2mkPtXLM4hsCGo+TN1EIeBKNDA48RnjCACLB3yPhXDSGXM8xSku6HgYEDocvwixPM+
oENKGPzLxf8A9Y3hnttUq0ztH1r1E/ZPP6xJbCFoi1+FD+nW2cRMQz/W3xVHdOUWny/CpLswS9bf
0qzf908vG0rmLgUhq0tkAvHkmUPjpvILHuuBmuntQRpgmhMYZOaZDy8hJdNJPwpha3lkApfFbPks
QZdgzNKA4ZUjn5SEUhbO5m5VrAw8sRyvFQjE5j140bqb4OMcQOTrSxoESSD64vHaq9Cqc4uj0NwM
Lvetpy0DhVh2x2eh/QivsngahHrGh2NMwp8+3ZnaTImmVv97aydThp3oxHyaTg5MtZrvZbdm0PLK
30XNEKR/biBwJOBrBWGmqgxQ8HD5Pkvfvk3vlfoGFf+5EQ2JoQUXvjznAFmyOA4okFG0gxrta/dw
GJQk1BlPtwARbBqwXRpQE2Al6ou93PLJ2Smk7gdFFaA45UXW59o9d1R1AXgPIBrVLxPjo99Q3kC1
1136PjxML5E585+u3bSWVbRLxPK3hxuNg6NBM3EvQQdAeqt15ECEVIrZPIzwLed9lH77CTISnv0t
R5LX/8S2xIAas+fXe+a60dMWG3lGUOMS3wnhz0gSOg9Koc9CDhhGQ9wztAuj6eyQzeU9AA5PTWQE
bFEYc9gvSmP0MrQZ4CpgcYDgLd/vR/fBDON3/OL2ZZYQrrow1MKGNmJr+PrSgcmfqVY4dcBOlMzu
/Fo6QHB86zn7Gw4KB984giYqqbrOCFrre7J5dbhAlYj+zo15JJwKRDwgSPFCGOiKA6Cij+4l1mdh
AbshfzlYgbayo2HlwyUK6d4oQfLYckp6LMyijlsDmv746TTzduViXqshn8/UTEuRPgSSVrwSw1qs
Bx4i9dBKA7LVgMcQC2/nKs+WTOqJV7hX4s4m5at/AF7f6ESCRn+Y8dClzit69tLc95H4Aqa7dypa
mUp7ODSGfTro3eijZFEemHmfBXM5UtxxpSSxW0Og5dVz79zC121uBfBnqUjRh7POCsCF56gEiATB
/XBJw4BvV7us+WF4UFSUW5vY9J1MQkk/OUpBX+xJzqWZCopunrXbdYY4K6uiPKGAt6gR7aUc0RWQ
YeSSLoVVJEUu9HZcLG919n0ZmI4+cEloPxvDhmGuPedYoqg6kQqe0y21OfD3wMybujNH3dThsR6p
qNxj1PoFGiHIGOHDsLfXW9Xl+AZ99F6psDjxIGNL/GcDgtZd+juBQtlY87CpL9fm51pERogWxgcs
oILVlotiggEKs7/maTyaunml6vA8zvZzhkId3GyAcY7ddML1zZdcwRTSpqCagDvcrqhzEGycgTgm
bZQZuvX816yY2CE2HpwcFDEjLsgWFGj1B6ZBDV8MM3rQ1TLfIAOpaRBIKqMg22RIiwAQBUA/opDY
gj2D8q1PpFFLurlCW6F4QKvav6AYag68vklAb0gsh54rSJuIETYG4vjtvFx4GNxs44IO1X66djU+
W4vWfNDb1T8KHE0kZOhqMaHyZb6hYWMjWYwN/iYZQVU6TjVbHVUiDYmhfHkMVH5H8udSwN0fePIU
XQoNXA3n2eKMbuAhMBoKuSsP0n7+NONJjxwapEAO5Zb81aVI2GzEUmTBUb5SXRcea6gbSh3XbCR4
F0JMie7+Zq2xEaJvo31pC8Ule+fQR9EjN+n3KvhbBbUqwX7CYqqqsbCTsm7pn+Z95TotXOt5lKwD
meVBYLl0iD99HWEIZdBsAoYGD6TWagj75ySqzLQG5VJVzLDrHiYhRhNgv6NLHI7UzQxw5iHcrjlu
XdB1EqLHBMX8FVW1Mp/9O30N0uqRwyszGdZH0DO10mHUHewB+vhH6pFSvfcjI/CJ7PSydF41Y6HL
pIkHpg1LoAbzXSQH+E6fpW1BVGVDc5gABGG5HTG2HgCGetcPfKlt4BsuWBum/LVN74xXuxlBUsra
gxi3YKb3Q76jLWBPRvDxnvPX+QPWWgL2sBvyE69sLL3W1xxlfNBSiF6ibhkn+RXCpzRQf2iCCXOU
7sMr+v7+ZDWUjTHJD8ww2wEwNAAYOBzEoqEvx7KuHZ0kdJS+2acu49jfbEphtCzT3R6qI+mAJ4K1
+nSKN5JCIlasMwOTNYSxJ7qd6/hcVpTiwlApjZ9SQcgLwIHxVnqm7528O3ttsVIuRWqx5c8ghH3t
bweYPmYdgbvZ3C9s2ZTBe5fH4gMwVpYlBXuveM/mm0Y8IiZcCL9x7BvLLmRekRLF4aEUDYYF7r9a
bT5GqLthEy8yQEE7I4T4c5dVFLdLd2nNnU39kqCWazy1PqE+qgbGUD9k9LGwa98+b6visSoxt0Dn
COCspAxRBznSA/SMqGmkQwWH6CJYbdgGNzGmzfcnVzwOCVCBSlMlrr4MtK1o7uHWLLE85sCVvbhd
IhArXxYdtbtV0K/A8hxFQiAZhwAOoOo93CAqwAvJ/MoEREos0XObrNKTSCOjstTe0lLJmEqZSinK
G4WKj+51jNeIeZTEpbzWAyG2kTuwg9hfdiB8MtiRo0C98Z3E+1adgq749Jm/LDEXBtDQKXa3wKIp
rQx2bUSeoq0yEp8e38SVTIxKnOvueOp4rJ8WAveZN0cYjp0dUNAf9tKgHz9mIn96ySDqZLGD9Qy/
aqjgcDobUwhcP59BvKbDJdDW8OGmFPNAZ+Y0uP9FgWknZ/Q1muWb14zAjJ8qBMv0qxFqL5UerSIe
SrLeEiF/CZqaD22ltKv3GXNy/wjqvgUy0yMwQUGXt1ZHjFSrRdDjdZjMn3BUOGo4l0XHJ8AJumj2
B0T2nPjS0XacSxrnE+tRAhNJKa/56vsrxELiSCTLujwCurrDLoX9i2sOw8jiOAYhG0BWMYPDkvTG
u3SvBmdWqgwyWSbQV+Fez96ibHqBV+cmgzu68iYVFR/dh/rBk98Dw/HSzAYALkw5y3n0k225OGja
pK1TUsQVogdiUkiThWhab9Eythl1kc4Ao3RmGeJHWcRXlU9SrAo+kXO+YUo7/GN0hR+K3vQ2kkXG
dEythETtuCBomF3xy4eI0T1yclWD+gDGSBTJB1YPa/9hQF7EHvf1F9U8ICjDLHG/x608HOHF8ArO
B5MlIv95gSnmpLJfJfOT6+9gClC234zRY+RR9QzljMbH5IBopAzQLyaC3lA/RN+5/mtNaEWONmgP
2umq0GBXqfqGaA4Z1tb3AzxcDJdjPAxZnkl+dX36h2DVgu3YXzDoNSDV9WzsNQtcaqn5KcIIEjI7
npNCay7Vem1jWmtJz5ZlxjJv3Agt7kP93JvphnM3bKXD4phXCoQtniPozGhlWC7nJlEaXLdXEkdC
0kvi++kkQMoszqwCTbjjfNu7QUkesxCrfrEwwBdnql9jHHhZp9uzRS6rXIkMz5aATdQSLiin6Ak1
JCu26Opf1nu8TaBMwXlDz7CxNTFvDPTw2RsltdYWKTx0XoDspceFgEmgNSrUkgcvdpCfysvv0bgG
iXWSKtAH9MTmmGpNz8eNKuuZEDkZEHgpr/3KUCvF4OnUvfwBKQHzl+5QGfVUaeVVw8E+lhg3d5Mk
crwC7SY2IkNikhZ5G5thkj5k1GA4ejB5ss0fy9ZNVdRYr3TaU3x/bV9H2LDhAIUxy3L/fPa4zf1n
pxtTmZH8yWe4JzechCeYLyIytlKZvDRM6ZPwRi2ltt2Cu2mtxZ9vjBAq/JqMVQ9VnBQuquMQUkkg
Upxsy8rzmWyJLB9K99muxzkWHsN6eHFL9/ia0Q7zbaG+A/wimjdASGhPiVe1QLBVtT9s63f/sJiX
RqjkXKnNEKOaTqTXEhZrqpafFA81AL7XcJF6ni6DrwG9Q0+no3kgoKQx11EBAgXQ3jrDInGnuIfm
St6JZH1DPER9UkGBEdyHpbuwk/IIkJZzVcUCmWdRK+XMUdqLtLTbxI+pP6KSoFGQ6esTMRx+3JsL
rEsRf68AH2fdYOc8ErwFOFdkkmygQwPn6RSNdVo94IrSavUOBseGP7WWQGBREnpl6VKFV0U3e8zl
pi8jfYRs8aQZxhnTFblkOCoYUonim64Ce/qQBDW9BVuA06HJTLUREOQQnwHuVoQZjpg++k95LOhu
niNLiyhCux7Z1aQ8w3/97/owSiH3R6FRa/KYIXPkmEgR1UnsdgIvE8g+v0NpELXvPsB0GFMw7pf4
5hphTP+6PzI9K1mSDAiITkuNt9dGulkC53tKjog+NJutQUSICUxRnjABE1HsUj9XXw5/FB9sSPWd
eSItfgV8wal65c45pNoAI/Isf4JU6aj/4+3fcOfhIp5PbjhktUgrYeV8xUACR5Jf43wNnz3L9mHU
VAWEM4zA/gqAKYVngFdHHicXK4wHLYKmAxBNdmZFmFsDrrjEh/QphfHqhwr9tK9eYpQFgRpMuaSg
BI5JWt0l6EuS+TK+Me8d05VK5K+ZhxkzLYpWthJVAtR1v+iCadiHPKtorje0qB28YFgR6ioMPSgN
CwBKrEVNaIldR16LbytvG3LzGTxdOM+EHdRkyKj4iTY6qK96k0rnfJhRrsYxspkLVaAic7kfoyP0
N+EGBnKrftwy+3TLQyH3LLQidj1wehGA5fI6fE6NirBQZf5h5Ssmt5TSudTYsxrh/3Dqs2PhQtPA
WllpsaCYjaw4xSn1TFAshfERhtCHZpjdrO+wVBIScM6Vm8IVQJqn59Wa8yWiYb/UYtaehrDo+UhH
iTtNut3TpaX6LbiWlXG8eDjJ1+hrWdIoJvCaAZMBm5cFvmP+Z8OSKg8UsKf4SbCiQ1lYsArvCRL3
p6UO5uqqLhwx5A4wfwSXEHymwP+dBp+4U20dC1AmlKFQQVCj1qEW1iPs/kgjA6hMOsNTbOspw2Oj
oZIviIifeHBZjZXS17JAHw95iEmhPXR3eZ1bwjjoqcbISaGKkIrS30lxamUpFEqZw4rEiDdW4sua
NhOWN12yUki7EA0HRe3Ctv7ezy9Q8NklVNRQCm1VKn1DFN42t2dyMYHW/sBl92QaPvsZcfrpbuuW
S/BUHTgYs+anmqaeXznWKQrt+AMoAzpZ3xzNUByx+mTbh7R80Jgweea8Z8FiA3DaRO0hUNdu+2xt
sPFzA3JADKk+pJ+vX7PlLfwFJiWOAcke6aiMzoj/Vnfkx02e91TO3P9eOGdIZ21wZIwK5XAPsrf5
FiOF7sj+hbqo95M9imboEy5FZbc2Qivs/E5FIPHjKuvaA8X7BV2tMK1IQordO/ME96ZKbtYDBm9n
J+e6nW6up/j2iBq/Yscp910lJWRLP8sK3EvVubuezGqeEsVbhH0GWbnfewBg/O2hRZ5u0WwpVrAN
0mF2CTpY3KdnU7n+PkIUeL6nn2Xx09FDd/X8S546IJcdwlT6CD9Kpw6Ex7FlqApwshNl/8QnC02q
lKbydBlSaVCBiTT7umxbpINp3Dev1ajF2Hlk581WETuBZbQZSB6AK5tsm7w1Vdmdod9lJJfR3e15
3mzWHP52gNP3DFNyVzaqMsJy1ZJyviVJVkM7b0Fsx3UG4ELVBaJGO3GX8CsbD6u20yB5ZIbz3YkQ
asuiJmqwXiQ+vUu1L9iQ5yU8mreImfwOS2pu419FG0NotBKk4drkeGlVE2MqpCr15IPB1N68zPMB
HOb500O8EEQ5xaezrgiqc4vpioZQVg42K+0ISdPRXbE0wZgWa6KB3cp2+wTiaJ9IDRod88d8oXmb
EK6rXmdg/QW8BQ+5Nroj6aIP5fnvSqqO9rmhA8Y7jJdogsz+LNmSTVe4tFSMmbjp2fRI2zmlQ7mw
eRF1Xf7tIkEdDbUFbSqeR2w+ySguVOZ/debK2KO79NDtxbXDYcL3wUgo/oHBsDet4EjGWmW81kfi
SaqLhfNEwtv+/iAO1LKciDKTdmcSbqRSHTr0JoEBRbmA1uzswhJuxlxQKdSH0/lOtms43SWoil0n
pJN0e4utFYQ+Kmt8OiU3mMwWOK5FpeMl4omHcTTrR3kRuskHQHg3EZ1pcXHJrGpiwIkqK82hdoWO
tORMKnVrqTJvIsWM5Yieux6jWg5atxXrG8LwJIYQE9aPgAVxnFTN7Rr4jEAY1IqI5njgCScovP3Z
5URo5XgsX+WSJmVD0bEI9W1QZ8aWzXoHG7cWmpJ6pN4yIt18tyLi6WA6uQ/b/nJ7/tKuqgPeDPJ4
Z8aw4zJIqPfv4oRut9tP8TYoslkPxG7vAxuI9p1Xt2BpypGswjHz44Zh4nkFteHe9IgWHZkfM1TP
XISosrN4Cmeurb7orozjamJUSLRfyfZNSFisUGMw/YQaZQXUyXkvhUd21ZP6rudh5q28HVOSO4c+
aE7U3asyjG9Enm4x/Hzks3ptXhKIa4K7QwcWunewR6LWCUJTpF5AL316qryuEn5r9IO88/TXcfY0
mWhk+XNCSP2qgHi2lRc6h6SbzD+i/b+0mFwyhpJn9DfYPKgRV2WIxUzX/IRMmHGo/cR6z0LGT7MT
f0xDmRwsJ2AA5PHl7mA46L0Bp+L5ZBZeWWH/Kozw1KBZKGCsQQ4wWG7qFuRpmdhpWO5ByZfk5yWT
d8oAxVTamnLmwBWUB+bQht4AxG1wJ72TvtsbtT6W5gfrtnvPwYqiRvjGpnusfxe9CweUvwXAzN92
rIcMm3kCmpeCgqQKoMXC9coMq+eLSqCYUdWYimLeYJuMynz1a1Vo99LxU84FXZAvJR4XK5F/RlRT
KUFthdiJtuFXDerRzK+k6LexvFvYzn8BhR8DdpCpcLHEiu8tKnKMqn36vXqAimEWIqTzv18B0BZJ
6lrvnXo4h677HrRaNqs5HZC8NVd4OfO3HV4kM8bFRrEJ6YL8IP0Ze6LYS03M/Mf6dzeKdWW7hztq
fxNcv2CbLbtzg5zdEV2/rJugF8fqcrc8nCm8vK2mqjSX9Pz3moCENXYVo6v2M1osGj6BGamlXDha
uki1pNgeobfq+Shh5o4HN19lN3C/G4sI2DiUDg9bhxtvxMPgw8Gfn9svyqSErfELtLp96LPV5ADL
7YNyWs1m83LKhxeW0cC0XPiQ9hEazwpIHrxcT6l2qGx5Duhqnil7dIieLn7a1KMvQxm/zaCVFGYA
hYYM04Yg6K/ICj61Hoie9a+cUThSLjGyeT9YbM4065r6MLpFntzQSVm1qb3+e6DO079mXO6xkx/q
hrKoBVDFT/DxrGmatwrAr+/dEPaSbw9cqvwCfTQ37iE8nGUI2HmCG3Vx2MJR77q8v2nfOgLskvJs
xRk5V1EU07yGXyycyZFKJOVo/TofDdSiumEYqI6ilPU8SntCWjWdWcdBPVIO0EhOTXGrYP8kVXcI
d/zxtMv6JLC73NzZ8EeQxwILW0kCEHre9sy5yr/zzyn3BS7xRWQ/lG63RWZbbtTiubSpYZ/jA+It
Cc1GEmG633INzaX56loMgLsTMMe0yRpGsFQw7WXiALsauhBEFzWuZy2rh5sX3qFkGHoVXH5Na7hT
qIIoB5QpR3Z2E6n0ysEXrqLM6U6MMNhNLi+WJbX16g5qpa0kPVTiSJ2XgZjsCmBJ4ypJ7ELDPzNh
J2ZCKuEpIpulO086JvTl5KzhiKQLwQS+7YTL0tmm9PK/WC1nj0lB1rv5SwSKhkcngiQbufT8Hdmr
6OpIw0jJGgYrEkJmcXfqdEI70Jos2MNm7SqGZBxKhJc7Wzaubk95RWlmwsE0V8xjJnZicY0Gr39m
cYTM8AGGLduUNnlXYScf64Lmt/pnMA4KvU9cDdBu4khcx4neTCXtK51BkaNl9XyEFrOgqKQKjaUA
JUsj1Am5mIacycE11UgOBN2PUfr4lx27nWaEVfrriMY5+1b6kv7rEQ3juFxkUKY9h3gQQ6CXvkHW
YVEC2qiPdjdBjzxJQ112JxI5RWU2o/3d5U4soyCJ9g9iqVSChx50A34v0vnCNP3VRk2SGmaNiIAH
Pg4CrGCJ+lPzL8OPbEnZFbcoohITrlLk263qAQBg+ioaUiGo0l+0eySQ4NFRP9SepsTcA9PGjk9H
XD9/PjoS6sCN1vwvUAkgw7+Y5FfxzPQTTFOhm0GM1ir3yhC+ubdrPs8HelX80hX4kapSZw8TJvOw
bMl4W/xDHaY7mKM/+cZJ9JHP39J+if1aLQMxlqJskhUSsqYjM02Op9xNjMzD5wm1jOiVVIoaiY8m
ZtAxVgB14/ja9DYhIYEYP+gZI2MnZoDnsPjVrvPWR4v8M+qW/8AO1fNG4lR+WjnXGsCr4ev4lgQS
Rk4C1zSQAMTzqwVZi3Yl0Lc3o+PRhlhSVr67pjIcixEdD6X8ojtQcDRjUuf2PvcTWvcSfecpLzXP
z9RVAJArJ87+fLMymtNs+0MTwH3Z0WLvfsbjVOUITmu2Ras7oOlQysjopg0xjw++hu91LWt6/U6D
Y14nn1JaAy+5csnUl2Wz/VL95TFdjtptfPE5EAxNCSBbE0Ew99HMFearknBpXT1bn4iLoroG93+n
J4tF3nnf/EHeFyFq+YZtupR7tcSIdt/6gaepNYTtZXSgeG9lR5LWIWbYMktwXENjPF04131d/4Qt
p9+CyiFP3+FYMKxldC51bJXupzvYm+fKk+w2pDnD2PHB6j7cocCUfFcJj17Rb9sHdh2ZFT+TUN8c
flI9NxuFwxMH/smk+lv0eXBxhDtKJPnlCgYl4Z0NShgbxJQXa7/BkC4DpBe2ejLHPl0ZdY8Naqdd
SZ/ZgU2tXFI4MiovD6Ux8sZ6HiGlRcDgCsD8reY8cBHulBbjMQvKLyRCczvFzlVrBPHLIt4eT4I/
b5hCco4dpzEsvVo8suTMOJLJ1YSjnppi/F6md/g9P+AFDu7eYRrfmsPgCfHN7c7KfFFKK37y13SO
GukRCniGx4Y3sC5KPXXd5xt8IzqSfCiT57/xPjm7/RPoEH5iMh2ob9jOlQ0uHa5dxnd39MT+1NQi
GsdXC8EJuSX7EcxFe//Qgl7IrTkWRRb77MsrLxgtT/NyxM7S8Wgexiuu4vIRgl4ZnD2jTpbnr6pP
izRgZIyW6IzCiqaNjxrWUiG8kO/ukG/oxwzF1gA9nKBM6tgoXPwEwx5hb5Qdg7kArNXAgpo6hEeZ
pGsBaogpVEO0AddnPBlxdmcYFzwyq4VT26hjVyXzvQBK7sxTU3FeuL9wi0etF3QIz0j/hp7jwTKp
SSSePwtyZlap7g3+2wdsqnEsMYWzuZ/tNuG68iwitsWeRJguBzOM0OF+tNIpaQmkvwURuBFVD56V
fOQ+a2+TPKnGyyhJwfaSthELPgV0USrwOK1RKAwyKCef2Zf54SlxCBgpneSDYjU+vtEclQQRLHS9
xuk9fPy4aY+VeAqlIiFNvW+dPZ2pBIryszOrtFQRa4A+8Q6TYGO+9BK52Ca4UoenrTfSOD+fg6wH
Ty3XNygvUgtBbjahaioV5jkwK4UWczVGXHxMCF88IwYuyqtRR7ZNXRVrFSSYHlgPwcEMkFlmD93h
kY4QJSP37QwJjptcnKhnYzDL1PTqUwmzDV+eV5AKUUImFex0+OWrhvbpKI/Gu+jreag5VA4Fbx/I
oxvwAIJ+13SF8titmfAFUcv7acS11Z02aOTI40qztipJt8M/QBH+ZOiYkdm3z2922ceyiZay9J23
mUyoc1vbD2yvtFzndoACzhlf3hDyIxf5DA32+fpdEycAVLTflJaEbM2V63ZVbT6bAw04cUHSWjqK
HJU0Zg8fgsT8wrCPeK3+0dsfHchtSxoarTu3IP+OeeL914z1maYGkC/F0LME05zDdf9amrKgNxKO
TGPCCH++jk79fADVlsTqOvWWbCKhsIsZHW1qFU7qlRyeoepNrClCDHXcUkDb2CS2xFbxc9wgJT2o
VWbc3ISTqBrd3N+m3vXgSrreG2AtJFT4O1nJgww6reoY+AI9TEp7aC5Kg7IIQsrenCg+w0sNpOo/
egryVukUK3qLMXhkwBouHMyZPKQHNGaSsGFAhlWc2vce9r6LyP7X19xxr/SjaV3ttCBYoILwQ86i
wQRroLNfdQtM4S8bTmSvRJlxAvn/bHGgIG7GB4zyu/F6hm3GuzmOj/mKg8rSl6ZgU+DLMvfYtWIj
44x3cGDwAU72Pw2lqOnPZd9vwGfYqVnHb33cvOW/DgIXTRy+0Z1XPQDqZc0zd4BPN3u1qINVYAI+
y6To/r66NKjNXbACWHuSb+g69Q//OisxeDHOCdi6Frliy9qc3mYmYi6LTJFmM+imsU12b6JxoKT1
p/73/1fozVAJ6rFzVFrHymATaa7qh3W0wjCElbtaCtxrryHk3+kH9KyDIy8pFgkwon5Qqy3dc16D
KBjXuge3t9KcBKhxSdqAWcu5CH1lBKMKQ+GDa3c1sN1RI1Gyw7z3s9MIXwk6EJSSGoEXUYplzc0O
L25W9bUiZEX+lrbhtxFHuVgjQ0h2uxRoYBuumpgAnEiRXXgvhsVU0Iry7FOCQhGxsip2qD+8z3Pb
yfBdD7sSrS2HdXffzAFyhg56PU4Qm0HjIBsClo/GsQ/WALpu7c8DRFM9dQA9R0TS/elMh5Xv//z7
MhA1eJTJThMm6vv/TP4MLZOsvc2l1QY9eMH/y+ynHSg+eAmCz2QIj4eSwYXviICxcll+IpJw9x1m
KjKiHUxqhpVgaD85Lm8VTUhH9f1EJ+pTZ6qPi9L/2TFJKEIg5KViljciU7UJqPCDXzmQ9kbMWjfs
TbFmO1B/00eLBaXGC19EyV0ChcYYgLzP8BUg25Jn7XC2sjovp3W8SvrjyWaegMT8lPQqJilXzG/D
q9tYgm7vciV4zfo9Ha9GVw02z25Zd21f5MoPZTIAwsqqVv8SlYvcMnwrkofhT3VTgWsx9RoiEc9W
96i6Sma/e96KYrWzzsV041yjR620CGjDrhEaD3Xox77yweRaShN1j4Wr09TjUHB3rd8w3kot+bAy
euv96TV+tIqc/75xCD7oIjQj/OJ9962tvhGSdP3Rt9SMmBtc5tIFCoOinAujJhFX0mbF1foGw1bP
zJqMDf2HairujxwdX7xOXKEJCIowDsfWm4Zrghy4s7ymmo/gChGBvnTCuIaPUDnJ68pWXvpy11T6
Q2+wUy+A1MjukfyK82mp5EFg5tlNJq/qa2ZVNfr4QInTeiVBqhW7lj8cSk43Hg5Ir2XddpaMVSYW
yY+FJ16ytUfcRc2gHoriYEb6tWfdJe31NCPv+xyRLwvcphzLx7H/lFMkKfh5ToNT3QW8R9kD5/Vs
ibwfYRK6oJC7a1ITHeWKSV4qoFl9g2/DRIjcVCtd6CFnijdk6axKxRjo8GAz8Fp2XmDTE0QvHPnA
EA8US97kmreohl1oO5KcEIrfiYgBllXRHlhZC4+CbEVe9ZtzU5hNeG1SyXnOFzHN4ede4OWXx74t
5LM91VffPgGOZQgQGCZFHSdvk2sH8irqSDpVhO7ETjsKRHZatKQbtG46sTSNukfbPJelhspL1x9F
Jaky1gwvbSVH8XyYI94q53UsUTpGqAVrDsBTgxn7CNsnk76nTWwAitx9cHRexwGq3Wl1O835s+3q
TJlC7bf+ecsp+/j7PkxFNXgg5/q8DNx1W1nExCahr7n87LR9e4Hy+I2ZcTJvKVCgvyv32eVKkpGd
FYDf7M5rClJo1t5Wsbp9bb3Y2PqK0XGpLtW0qsIPO9dieajCwK2xKX4FkXRrNuhn0xVpi22qTcph
dwhvB4ANNjdvO1JJgpykcE3YO+kDq7aeYh7Z3luU4w8qEaOSFyPJaSuB0oqQRQ4TW/fmgl/4h2zj
UHIYG93rSZ7JzSwkjpPZsDuD5Yj/U7JEa+Lpuix9PQIeccdVQvYbrMBAIj10adY+ml7o2scfYJjk
9N1IJb08p0aHLrfFRV6h0NSSEhI30l+jRcf/n/0fPi7uYNrnJTKxC50M1lN24wf9rFUznRT+2xCo
XdTnhkPBwQKeDBFFge2yqeqdjE4FcmtrNJeWeQHfeqcsLVw3tCKDYnzGyoPaxP1d83q78jIei4sX
zHHfojU7qMCbokt6+LVOT+NahOiEcHFlk4mxSOaVasgd1qbakdnSrNc3RP4vz7JLSTY3RhJs5lej
XIsTg9zYju13IbkPMokirFrhpA4hR/aojzGVKs8EDP+UIBChh/dAZrwhestm8HGR5w22GVrIsxq4
EA40swrh3cPcEeWFUd6xUUR2ib+QaBvWlxq+07RdfsSblZnHYBMxLDejqUV/IY77tfXJPvNxw/Wh
lH7c8jNA+g7+1kcjFlcIFLngTqahD5QCaemFDb+obNLnC5uDOg8ws2MceXBAjKS8Et1sb8228bBu
s5En+MMRWKxwcDBMAH5zBxfYJodIIXJZQWaNqsrNUEW1uYzzaoADrNAFQT7fxcYE1IpiaCW1My18
QNruX3bLDVG8E7KHuD+7q/NBgSmSu0HiS8pd/TUMg5zyP8ie/h5xZXgWaro10KJPPZno4vbp6ick
AtZIDy+0ID5HD1qvmYcu8N77lXz/XyW6PkkjHwnszq8zCnQB4SDZ5oTih3zMCOF7MPMcAodhU6Ng
Wo4SXc6k5ouMxWHw9lLZwGeTZunZhAwaeZq7cj9Kg6//+bOOt9prrelgKulJK4o9ICiL4eW720Q2
alZGfkfH9sHOeC97Yaqrzro4+CkKOAjKHwFXJsPW370WsJPv7oeMP2ZSlv6InycjgEZCARx7EPCg
JFAFoXZr+K+fVzrwni0xNLy+WAlbej1kyWNR/PKpUhBlSEhUvHnv60mf8ClezLPAcGy5xuH6su/8
3QsDWgUv+oFtCwP1Gpqz5S1jT9gbQbGVio/cV/zboBpTfzw1IoeCB0BJ9DAIGZKQPPuFvtZHwMNG
y5ID5YinVknNvKg0asWuixC7GZDmPMjxwzuJ0sfIyqYqsTUnpe6jkW4TmRKHWbxQFyKyaDVTB6Mx
CENmn0IPJ6HAbg0ZdhFXZ7fPRZ6KhSMAPiKxC9OEI/HkGgJ89WPKvaMmQY19cPqlPZJqA2QtZ6Ip
LS7Y7XQvoQoxFZoynMQxH88BBDUnafaZyOmH+Wjz+ftOy/37WPj96YAGJdvxSBvFyqt+eafA0mnN
g7Rlg3gtTEdno7LtcAUTlMhpUNVKoC1DokFsWmW74pwoiOIUbSwG88h6gL02fqICiG7dQn+lyrsT
n+J7P6VQ8JbD4ywr6jAjItLehdLgRh/Rd9hyyGGxflJWkWx1jHYpe78Af9x33jyzErjTG89VNBfL
FV4w4Ot2Bwqw/5QYhnEJ1WwV1Y88nCImo6KZh8y3NPaxe5sDNOBWgMl2aQBtOfRIAdRSfXO6pFIt
fuu+b3W2WhzNIQon8ACrW/Lsj1tfJvNhQ8ia3SUjb+oMRYXVfiNsjQ2Ff6hELR1aj01B2bfG1rfC
SCyfIcsPCuJaPcqDKhST3/UFly/6PVkWBErzdAI+Updr45Z4ScFbUtaHRN5AFPKxy5IT17dYFthZ
3m1/vmSuRQrft1sPvrJD09VFNCc+AaaOt/3o6og19FP2q8ni1KdR75RL5c3HwtoC0rhYV5XTQPXp
K7lM6G29ElcaoyalRNAnPFimqDivdXiNtFixW3XJ4RiZ51PO1cx+0EH60TRTkqANLHv4kZy4NfPt
GFrJRkYUFs7ehjTY+RbR/nBpyAQZz0oJwz/Uvtt6UVThzVnWrm95QM9ruTyv+AQkmCekEPhRKSDR
xe8s9fCH3Rs+gBAbrjjw3Lcmoy6JKd9u6O3HUXqzwV7zD5CAe4g5LZuCok2VlbtnpsfISdV/H58d
NnXPE06d3YuEh9u1HYYj/P1O2tYP9WVNWiJUZs0wpbidJlJQgHWVUdAIfp8dmrwMU75AoZv9pVBt
jmJdFSB9UEvPdw+CGxWr+hcHQw31bpYQ+Pskq2IN4qcSbgRuji0rSZeMqghRVIKQOPgM28x0e9Lj
4J1hg4F/dFfTym2RYicBjfGH4hqL6DuwAESIcqczKjHNF2TLDmKOLGJo4uG4L9LMpBjezI4snZlU
axsUOzjF38gwO6LrWEmvXKVYUydGuTW3GDnPsyDdIfVIRXcnvhht6zlDM0mhRaEeo0eDihyvEevc
8jiUWQz2+8/MG65FHMZCKyD4/tBrITv1K3YbYiN/HXgzt3UCw6UFrjxtaum9CWIGsbFATnMiAPdc
1cc9F6tuBBxB6YBbIq1M/e/jgBHiNrWAAZ7FU/5xdzMV6TC1EwNusnR0DlED3Ugxh5wCYagInGO2
40CxzjHCDwQBWPdAgDkDKVSrov30SpbDsDR7AQyg2doRcB0ZBPjOKq3Y9P3QGREV1czBjofxBSdJ
L9ZDEpRwmzkqvc0e7CZA4rl1OZk5UwoGhdzJbXqB23C62J7wmkyX91c5+NEryafXXW7QeN/k775r
F3FqSRKjk8StdRAjkIRl8M/Qf7/+DE0IVnw4oOtzTwjzOUwxERnU+NNU7Fn5LMeHom8SZ01DSprm
VxHFUGXS7AT+c4JFJ7ZL6Oxaf8soxGqOPK2I6Rp7MRW8KtmK1nUh80cAaDtZHflfuHdKYDAwNW87
JsTAQay3cCXhR15XAmcFx9hKdwTCZccv6kYLG+y6iWGGys23DoN4n3gLqoQdbrkOODvKFz3F2ppB
lzOLZplLotxVXPwlnMXNiVCgPjfpTQUY5ffgdtov6dj6GQ0RJS4H6xSm/zGMs81zjyBa127ZnLjG
HjJtwDn06VKBUXmxgwJhL3Q7xF9UpKDEuLOHW/3FtUpfZNa/luNp6wQ1lnWNjNta/2vQ7DbCq67Z
vfIxT3geG2jvY9d8Z4E7wNrCF48Jc1gCQ7UHNBCJ176dSfoyDO67zoNJdX1G//CMbpcpLb+jgG4l
tUXGpvSPNxJ7gpsuYx6fxpbIAAxLaW9P0afzFzFOb0QyBE7uawBV73nbzYga9Fktmt4HcgLBrlYO
NSyqDETME33bI35lv5j6naIjwlCk0mky/BZY1+nEba6vHQyeSASxvvS28uf7ezR5Vor/2tl4N3JI
ZRvy9s2bLDyGsf6hjuY0FIurIAz+Xbn0eZUeKJSXNbvp8S6yByh9mISU8hEklsmco3PhvaaQUdrE
Ut73WhS59w+nST+gXADsQ9EhZZzbjwuS0fwVeKk5vCoM6WR+wFFNeHGyxndUOwu+LZtq/b+XnmFL
iuv/gwGqXltQnk6m7oWpE8EGrXi5qbfQXovc1Gr1UkC/lKz5mK08fEwLVG91JbeeJeWNUvgA30VP
kmr+h/TaMQjPmGhIg0mMS10bNsdyN+rdJSJdB5PRAcPW64LP0uO1DcidTaU70QhxfN0q3NPFivBE
KQZSEGjHAtduer1dZ22T1IKCFEbuneQVirCoHfEQB3aai+tdGCdNsoFjZ6/oBB4GLOpUZUKf2ZXR
9pKwgD0NTwUVQ/Xq0qZu2p1Qg3ulywJWQkttI4I1clELT50UGIBQAenPGTI6JlRJcAhOpxQ0K1cY
Q8MYFq//9pV9loL7cG08epg1dJCngbzSj5A5k5c9OL8imynoTzB6u/4kLSEHpyr6VIExeAz3ezc4
X4vbc6U0xSPm894Jewth+w5u7Ojkw6GehokivJpWCKH4tpEKpRNeN+11/jM2EshrOzfVT6KIDOiS
swdwJDieeHqg1p3pfaq9CTPiwYU9nfSEyNduCa4Pyq/OJeY3O6y8RzDiPqMQgVXiWKXQTGPLMTkm
r78F5azZT5fH9hIm5AVPoIWmohy24OIurzQr5y2hH2dkCDt0/vAqLYhpaNu7i+Fvk5PHZk3E7Mxx
r9olIjTv4XxS/hI71nTY4Yu/ABOHsJ+Zh+LQ67A94xZ7wcQMW9OV4lNcSJV/czzJlHT0cVXAbKKT
2G/69ORpVbPuM3SKmppDn/8QAmUHHsFPuDb9Utvw/W0o3e5iQe+19UI4PucaU0c9S9vMEK7FYlA3
roKdcyrWAaOGNR2rSDUeZljr86k/YE/VQLCVOlAgo/QGudA5vNbJA4bgUDduUNzSnqezanX2yhf6
y9XdlOo8P0BQDXHueYDUEXBzQyGxxH6FrvfMNFoefVppsYE0Oitp6EEl6vYaR5Ckim00s3kjee76
pDHUO+2cv/tznj79XM3Cm4xJGMDQm0h+k3PvI0q54J+YrnTCin3jVDt2jW4EbwcnGVL20DlsGWaV
UhFrAJ4QfWUiLoKZTLKElfG4ik0jsE0zNo9Zk+cjkAAc1GbCqFyG4sAbYrOEqIrV2LpoMrxlOa9p
mRyfIp3X3kAWTyEvztP6gVUB3VK4ElU8f6kibm7H2yBo9r7fdcNdXkS2O9UpJVZgk64X/9/HDuq9
mVit4Wgtxx08mt4oilB98z44S95YhC67y13g2CxQB26sn39DGzSAI+AImEg8c0xFlYdWt9UXEsdO
3XN8lpdOR9k08kmo5/wFaCUgBIgE3bNoE1by486gOZisb6q8xRpUkb9TEuKiwQTICYy/zJHBzvDw
d9XPh76bG1Md6AO8ZvGkObgq6TGublyloAYTWnm6hY8p2CodftVtU8zymvzFfRFbd/pO9NuQ8JIJ
GUhMIsYi4K6J5UefO9Y3oXJE692LqYgTgSQPPi0tK8aPPflec7cuaDOydMjFl7xOlkMrUYGB2s2G
OGLsffx4RQh8YusrUYF375XrUxz4AAliZRagVhHYOHoZx0cEZRzw80Ab3TBfbiPii3R8Ak+Ej3x4
ukJbUtVOWQvG77yX3FIKGLXdxtvmTJKX3f0fBXzmLh0umMwW/1yB8QvkVbDATHz3wYLazytfSfuV
HthYeG0Su5hwjQuxi5OIj2T1lMihdzDLLRXaemQEpW2zRGGQOFIaJKvbBxqzkAXBdMgpChMhi/ZD
eIECoibtbPomOT6ycveN4MovV9LF1EWY3KEkzYgdxwptAwJr4TCEKvy0iwA5jD5ySCJScbJVpQg1
ONMhPxzmpwTNgXuQ1662gmYLL8zF7lkg91v0ErkQ834/29BIodfkAMEhK4SIlZ9QHNxPSvG/uspN
k3kvhXEiRb4h7IWhj2c5F17v2UvVyI5mfHLHxdLi2TvnrjmUm+U9LS9z29qkjLGF9DRvtsKFTxR7
VPBS5jNRwQqeGzuQUcUOPyjj+CqYLnwiYZS9ztCeMjBJUVfwAgpxde8Oz9QMTCdYF8ZqCKZ3QtyA
Y1AM3tsIVhUmsyt58hre732GAxO4obVvIHLhLrIeQ6oE6bYs4r/7dYNIpiSMLYgI4WI5YcC2sXKw
PLzuU994EiMnt6A6lFZxAW1SoJzbbzOkPZOZde1blv3Ze/V6G8Di7WPrUD+nGPMMHDibLH3uzoPF
lLidJwf2zJTkaPEJZUo59jWDACbBfMbm7NHEU103G8F5KADHk9qOuqi/OoX4Gx8206co8zNEEySp
BDKwriG+L04n2FWP/oqJjR3r4esjdq5R5xaKUdLgyrkOoHnjO9dR+Ats0gM7dS74yE1Sy+RyfrJ7
CHCXJXkyA4ix2YfrpOA2P8ecUyl6CbNTqHOxEHLQMowUzEpV7d83ESJiiy8wi0VHNq/81Ga7R5c9
QXSOQ7v5FLgWOA3XqX7NYZHSA61zGjGvxyPCWWodkCZJAeu4NGqxOIMrnWNN/us5Lf3y953Zkzxi
QJqi6ga9/FWuBFTYX9NLNyyykhssw/y5n2cn8BA0B4NbyVuHz10+NhPTZl3LUFEV8YX98HIauQP+
bKvWFcNAW/4xOR90IC9Ng/ydXgXNoHb+OtUnZ6+YLYzTRgq6KYV6q11zGKhywxunZnx8Mh0Hv+VF
bdmrJYLwhm+Ox1vhl4vFftmaYUtq6H9OIwmig+XTsISRPo2D1WpJagQWArWbHC2Isf4fZmkhyjli
36vfEmb0LXQ8X6IO5EQxLC4V4hNVMr7beYfHtLceJIU8oKunQHPTGKVuNzgGc4TmEnPNFwQwfIoW
eQSZfbgfq+fBjUj9zCJoy4V9SRYkjkiwrjL9UuIWLMarAMKJsKO4MO2nBBX9XLYSZeA6JkN9NimY
UZ9noGIdNTfdG/ayXNGOMb94JY84r7P6WYXm1EtAY2B5tdBu1SIhbjdxEFOToVe26YCUqNnW5u+E
E5jPojHLjoFDPijP3TpAFB7+oihXVcFuMTZoneEfvBYI3tryX9BR4MGr4clqeeVzfa0SrJXwtf5E
by83ZZ1DrPiHrIx1s/C6InXc0st7sxMzdmqj0+t+9ImLvzLFrWzN/ToAa5kOOuWQQmHbdeb8tftN
MyQQB9vUaKnTTEBN+O5aCtX5gF2fHUBiQyZUW78Z7EJVAOYmSIOULxkFeTszZyqwWGI2aGb5/Las
lcuni5Vc/VTZ5ePX8H+JEgwXSEWrse9mtt9NFXaZEYD3w/tC51qhDXCcURS88cvcByju/jHBr1bp
gSTzK1p6h7hXzEE0/lrxvLBiDjLSPtfX3m9aFGxWCaBI/MsqXKqqgAXqvIGfYAj23oLcMGOZr1pY
4HS7T+6rwJeGG+RunbQjVBRszcQV+sSKDCXXeTkK35X+X/jlICavwlg6iZouhSeXRYpereBgGag6
8OIstRWXNBqrECABhL5EwNcX+w7WXHd+vuew79YWY1ONCr1kJdrF/bVTbztN6HLDXzpeU4TP6+yG
nu5JkWHJSdoBfmthoum1KEpZXjzcDl98ier72PqjktagcUcmYzWtE3/MZFmYJ1pLBTq+I53FEjpm
xWx/kT99/vwYURM7A05Wyyd/66dQsgj2r5065+2bq59CjQDSDdzQw4NnUagfxqu0aWwVosAGYugF
kXAJ/WUgm8+j60510RPFo6rh52+Ut0foPDAkJl7Azp0KKTij2SgY0eZIXm8DW+5Ke4K0gFTxDNQr
mz9E6hp1oAad8of3rFN1zHagEhpbKQKHzSpxBaxQtqpYtDqFOqH9e+FkKyJH8qwjMzb0oze3PhiW
OktKBvMlSmONk+MO+EAiON2CAWXFEcWlisx0MB2fjkQvWbHfrh2TZffPQqhZUUGpqHBts1JZBXW6
0+FZ76QtanREP5+aNUZPafpbMmLsOWxO4TbsEzhYu5ddWCVidrojIKu20CnJFaQ9wrNjJW721Rss
Xv2gVZWwXlsYTht8dyR2Lmdb2k2RtQ1CB1VIQIn1cVX8KTqi+p8hC7Q/DsiJxKWn6PXkSmGGrucT
u85cPv6ANNwSnqQ5ZhuGQFN/+XmRgNC1atmzAMqSbMGCmyUFI9Lv+ih8QdBvKTWeBYfxkR6KM4Bk
Xur9NJ0yYv8PyWPxUO2a4L3ayue6auuWxFEP+4xhFuez0nMpno6OdPBFL/VVv7X1elTjez90b2W+
c6JtPlrLUyg3h8AWGijSbfxga9HRWvyYRuT+pal03acO0Mw6WpS9VTff4arlTHvN1SbWhFwKJPSH
CXb3bz6ZuOlchFh4YXaniUkEtJ/GXgz9LvVCCxS27I2Iyj1iUENY2P+SLzNi7IXTDhHU8Y1BL4K8
o8IfnN0gv3iiYjjuSMt4U8FMAUxUyHGoT4953hjsUPUAgJ18OYZu8SkmlSNWaW4ZAdtA4hIo3ayN
iuQDH7pqEE57AGEHu7/ben7VyC73VCbXClPuyBO3QhKeB9FNkxmTjznMve0HK2szdEmeuLhGjzJb
53vJZnY5qbGFNRD7PcvbT6voO8Xr8Tyq0r+8hsU/4CwuP2uBrm0GtfNKPEp86p+fsg7vQ7hieGkW
7OUo15x4EE2Q1Pt9zF3tnQTtxnOTGXSOQvrGtkjgpDvjJV1lpDn6oHUPmcb+aPAaZ5rSZGxArRRC
jOs3FmAuRwt9SBfsGhe15jQkeFMbv8H7rqGVy37PQlV6EJKLjNH1becbInuKwdIzVzewNZhmeCXi
CgP1Mgx3GbwNmK1XFBVZ35C62glNWXNmoNrCJOr9q7Upn0zJVfFFj86V3bEYGD6qfz06hd1yXb1P
lrXbTDic8LH/ks4/beBzARYB6lhsAgkuZ3qpKbtvbp/DcSzZ6RUgTQZmzzKDncjS3SxNj1fxE9xZ
BcLaKHXIGok7Jrr1EDWCkTj8lkuYpRarPJ1KF0hBu74R8Iv3TxkXLQ+syk3FiQFYeLBsU8u8Y9xK
y8YM40WKQPXNPCW0nBtAsYinEntZsgTKk6KIAp4jhOWatl8NwfIG8rOpdFWRDPZp8EtW2uMosSiS
7ipdXGJf3norWCgB6dijm8tBY9Z/6tMcN7uZCGk6BomvLmFCKLwmJ41siSBYQfj26JXCJGccJ+Zi
bAz1b55IjmNgaCAUCxC3wV1cedYqcYmzIEdE/FCn8BVfoApwbLAAE5gKZYT2ziCdyXmq75J7YYOn
/plhlPMcmD/N1DxiPfb3saWpsJZQ8F2iU1aNQKQpG+KrMl5NBA0bzbra12P3cyUoD3Zd7BuhOwbX
qHvoCVhLEnTtB/io3Cxmy9dRZuioVybvwFlgfExbq8QZ5TlMBMwNu1DGcOdugcRAY0fUKR1eV4SU
jCzYpiP3PWYigd8dBsgOZRc7J/YTtkWOsrgN+1QE8JQPR0sY3J1+6pDshU0w5FbSciJlt0LKc1BU
sDP/W3TylcexBi1S071EuDbfD804Mu620JhisQRG5/GiZJZ23VHhzTTB8O4nq6/yVhohwGFTpv9o
iZnpb0Q8klJYCtPVgJsSwh71jqGImPLtD3ZjLWArw/zO4WElfeHQrWpiicy4SWVPcARzDQxTGt/0
DMAX0nkA69+B2wsRjgDKNKJAyAg6Mf/Oo5ZjhCaICMgYZpn9uLEBy6fcP3TG7OBDNzVI6Mj2FgeT
z0RSmMxH4grE/myMqqkEFfBJ2T49fnW4mdmKRWfk42Ycyc+yEtzo72q1Iem+ZG23g05OLB+Ng1+u
VLpDtAORy2+FJt137KfzmqX/X757MFDFBhz3hO94BZrA/Jy0AF8aJUDhKuEb/tnqzTWMjtm072rX
BKqdg5yzxbppCxO0trmz4hz7TTDt8NZSeLHA7bodTNehwo1lpSEPzYTMnOWdjkvwT2A6Jd2WNicf
0rtN0ofhmE3Uj1z8ibiCUsfvOVLoR7ZYHQPPI1NfhCn0dG40ZlvUB+mpDldgQKkynCIOdhFxvGwj
K21B1fvqwJXZgstJcNgoAqf0DuoJzZDzeq8xqak8G40fqSStguUVFz8IU2etHM82e2v7sMzv7uq7
ArS0ht+3TZZ+m+Tsnbe9FmGe2sKKD/xow3AEl72dpasDW3AkJRiM+Jg/m6p3JoYan/QshAmmVvZW
yEyt2cmY7spxM1XZHM7opr3jGjOx5AWsZHl4+NjqST8M++7rjBK+TY7wSAO/CD+WiY/qlTkyN/d0
M1ihlEN1VhxK6+6hyFMY3L+Yz5Nj6IHj7A6cwRaHvBUfwMGQsx1M91Z6dmXyJDaTKa0gjoGM6LtY
h1cvcc6tw2M7iOyiXRnFcVxxN/GFIOxxoT7MZXCtwR8ivUmjGu32bTvAu1DS95UL2Qhubfh+XTBX
o09W6qHkq0xGJQ9OaGvbkYKYdW6TfKM1WC1C1dee7jsw+/LHQRwac4HqaS6SZ9bVAp66R/HLUvcc
U7JLitoGmXMk7EyGYCHN/9EUuVbp3G+q6Bd2yyjk+6G6UJZB4XFYCM4Ala2nuT8MehcK7TlSLzwD
z4pl0Buy+tVsH0LqCoQBYGqD/iIR6ASZTq7veKNbDYbAGmsjwdn3fg3x+3mZaN0a+YB8XyaqEwLp
wKADAN5OCgQhz2xT0VBrh0PQVj13hHz2+ib/YFHOk7J9MPZvD4mlyoIW90Atusu+D04LdbQcDJ7t
btjejSp3cFRaqPyuYzWx7HAU3pOA0Kg2WLjPuUY8W4yLE9UElf8xNsEHRwFdl1nemVE4QDIfzvtj
iT6XY1g5tT0sbH+E/thH+Xw6w35KMribm29ZRX7Jo7ytd5Z4rzPr4U82Bl+X2XNzSoZtjKl8fiSe
QzC0RaBtiHMmSwQ4kFokue0Og+2iZXrC8DZP69w6wa10eUzMN8SPYUaVBNanuw4xKXH/HOEGzOaS
z/u02CTQHOWP6ZXHEBk/4oS0+nqYOKgNMO9mVxlWNrizJMGELTzpow0QIRnp/oj43OMzsc9g0Iow
wKFNaPcW/R8ogKj1DawFFKmDO8sNnJQTqJC/W3lQGp8F6Cc5cBbgQyoqWX5IjGNgFvHsYmFy2LOa
axiNt8xKQxUCL7rzje3Rbisg5eFlZeFImfJ3Buj/wCJ2rZiglk6/e8czVmkBZmqCq1u7RUD4yqOC
ija7SSixzH3zuyWROrZo8ph6lZeTdgTkSqDWN+quHTMQKGck+Z/sBTwHzxnpTtUMUHemrPOrFxlF
OWyvlDkC0X4Dr5HCmTqEvg9ng+ux1E04ZiqIFWJaJ/AcHt6PLmmJvv0WV4UUdQX/7wqgr4glPZSF
Iq2etgTQVwFya8Ihz50NqqG6km4NyKQqDYs5UXmulN1m5GATXHblE0APlGezv0Feos0M2NhgOoN2
MDYUrqtBUIHgZVICFYnV86F2jZJ5tsiZGMrD00VjHv4E6IiYBzueqAbNieg14+jouZI9DnhTOYln
9xNDQqOj0UKBK0Rbc66YcGPYrz7zuTjpm5rHfqivPFjtWmKeWYCU+l1QnBmwASeNEWdWmCH3XYn+
VOyIcrb9KDOeIqF15JeWHQS5yqN+6CnAZfHq90AZ6/5Ll3kjiC/LnXTDKuhs7CkiE3Nx4HVXyyWr
0mbMfrekfQdSRQef5XntbxZ+dutACfp2QLA+Dgufs+7WSAsDJsSROh4kn23bekDCxK+NS549m0RD
6gG0TxQshxL6gAA9lgNDyL9E3tMsFIqthe8JW+jTf70AmQbTK0bXJbau2BVLr+PnYCHMIljzIMNV
pCEordjoj0NhXI11LzijWK4L+jDyWSSIqJBq4ZxxR+OSQkLLKYQVc0xnURU9B50OKW9mj4UMAzAh
p7cr9wvdOrjSgn7h06kO6U2/GlY5CDkwuobVYwyK0Mbw5Pxb4Up2aohu238/zFepPv1+LMbWDqCA
8E4JzXXu2H8dOLjCDfmFAte8L/KN5pG6cWGo7K7lx6bNISaxtkVsVmQTqbXp/BMbDahto4x8zCVQ
DYIg6VYRqQaxskqYeuZs1V7mazzV53kQkWJQTePmNp7cQzJIzMWv/gPhnc7HrFUTsm96Kd+mPMbT
xOCgitGO+MoR1o3hSQDApnIwzABb15SGyZ4VAesGKcZAwiLzNMFm9KG5ZToG6l0i0JnetawXW/YE
MRfpguFP/0/S2kUGfCzgK+JxUv0eBW/FW1NhvrEB1uQf6eEUAkoEUpoaZZwzS2ub/lPt7xTKrrBf
5KrlfKtP2Na22DlultDADq94OEcInnF+DpJXIJVZI5vuCCxLY1cZaTNW8ZQrjvRLi5G6kFfhdEBN
+DPFjrkfxi/I5O/K99zy3WIxVJdk4f2SzeWWhaseGWignB6zzDnndgZrhIyHPlyO6BwC7DUY2q5g
PGxBs5Hoitq2b+9W1+K4hc+zMwWY8i9z6MNuIyBevUNuxdoxs8vqbiB57e9fzBgXM9sBzo+B+MyP
jk3G6AtROjbfzCKhsN5uDWJhRX1p3ML9B/x/JX4N5yjMb2UFm5w9alaygqmUCL1VOIArXwNjCZk1
GLEA0JLOLMAcLvroNvGhlOmVT6dwwmDC9uwWURxWoYc2ZLMCvb9ua67na5BFGxH1SUZfCGuCr0kR
2zzn+++zvbYns48tGhQeOCtpAGGDvK+Fg9wi8AQm+LNKO8ly9Ya5a6mdg+wk4Bv1eCVLp7wEcCxT
vnumHy+0usYe2IUMno8O0+U3HPyHa3DNoUViVEfakWrZ8CACiLdbT3FCDurpxLg7j3uwIpC7ET8f
Z9JrOdufrFUG9iz/B05RYEh5pu90ze2EVSv2oVm0hAoehj/KDENnDF1dciuBeF6btxt71RLLEi+L
zcgQ0UaodvIXw5nwz85rHqoiET33vHQoy2QusxsLO5kyCs61V4wunBkj4JTml/CCP29/xlO0FEgN
DDQKW0DSspPbcBQxiTt/ffLvvcztxfmYrNiS27MRAfolXPA23zhkIURncAlcv/YMvSzbXVz/tFx4
ZVcuPEFL6mVE/iZ6LNHwaUrYMjbdCkiHvltDoOsn+WITvLjVAfKvna1ZPAqeOGXPHbqGQ3dIS5IC
oE+RZZxx7gXPoK+BnZbSn1RGmbtNAvnD97MltXoh0eTjprbZyRu2HkHFpH+f5DAscSp9VoKhXhlc
e7qqUyttt4HLxG1jVqrQLT0vljIfUtTsUszfRlEY9TLucQnuCM+0K3qLo2OD0mCCfjUsHzE6rnYG
nlCkupGWUZoybin4FZOm59D0hVazGHwtNX2H/DSuwBfxCn5VQC+F7/+a3x2LzVjD/crVvp4WWDuI
Wn0dXTKQCliRjHtBz7OrUQ+QvS0fN/MQnfdTkOoizEhVuhLBennJjU4ieZ6DGRxC2fFfLyqpeq6k
J18iZg85hlrvACcQy3Bo6rWeQ3LrifQxxujvLcdNtsPNXzcK2Bkq5bdF6Suh8QXIp/xo4dscwRjP
kEPmXTI7Rn3W0BA+Ri2Tbkbl0qSrmWJn8RF5M9hORmQLKsRgoW3OudcKfocvRERBidK+b4/DX9Qj
Rg+SxwUWhY1qK/LceoM9lC4ReduJK8Mu2l4cfF1RD58tGqc4KhYzTvE2XuzXv5leL8IfJbd3HV11
cIDm9j8o85BRee36E4OHslvIXS1IzA+YGcY3iYW8x6ZJpfvFMYZz51RV6F0sfk9g+UEJL0Eei2hc
zUOM35l7QUAyY43CWnbI5sj+/z/NK4mNq0m817WjLpfvXUZC8LOYCMU+IqCyagK/xuGh0jz1zRWu
S+jD5FCVXZaN0c56PrMGn6oo9qsqfKoHQYXgvb1pr/SPY5Gdsxdp999gV04my7JLo7xhointa2m2
pM9q+2B/zsfYE9d2ttV7C4EWp/ePVzuIVUv6Roog6TmdBN+FGkeoZ1xGNQzvrlkCbwY3L2IghQkp
x+lonuMM6h1V/k9bUYsZhgznW+RfIkaVM9d5F0o5hENtjge9J+lDkM5PM6EFLlZS2XXQb/wHMO40
p1fY3TQnCjJ/QBheQ+wxeCJdFsCEGS4DJsP09BaAiNLTA+1A81USRzKdeZlZ0kOAHsKIb9lDlPHJ
HYpGoyS8VSnWuBasd0AC7KravbF9f1N0AQaE260UaxWjgJA22u1dM5Gulnc9md6RNG4HsvlHtfkz
NmJOlUFaTGG/0CjZK+c7pJo9xZXB/SVhIdv6x3YCs/cnuIghiX3WaNMxfx72LbU46B9MZbvHrroZ
KFho4iKjzdxF3kL6QMGMfpiewz6XSL0QvPVEdV5JWdnv7L/BqBrhLt0ZHd5YgNdbc0DxrRNsY1kt
G1Zz46D/cRHYnz+cWh77lKyTD1JsFPWPSIG99OoYgF0dIpCuOWdMIbhq2yiu79WdSU63PH1KMCVG
+rLbYl7qCFGCrFYl7iEQlcLPJgw3fxpPdCu065xp1/HiCXPmhGRiT7GalUeVXza1vC7oZDYr4pr/
jnnuQqNnfAEclcb7UDFNHzmYBSrJMo8/UNJTyR1mJc1m4BM0//EGsje0/6rlF3ERiXndZvFPUVGF
ky1y3gO2D7MDUd+6FKIl1TDliELJuQQX9K2v/q7cHG+89F4rP3x9wag/9YbuYtNUIvupXJDQccc/
D8trFCfZtcLybOxEd9+/RdJLRMBybCvd/H5jhlOkBmCXFLvS/wguxnRYxAbqImpuaUKiVGh8z2vk
h1LHYePjwjbA6Yt24YzVjHo1VAjAFVNBvwiGLYLhsD2MypODftnonL9CibwPpwvsqFEoaHY9lWwQ
1TZF5h80CO/ks4G20ze4ZVQ2mNiA4+tmMswTPkpLNtyWlJnsQS97Jc44P9FzKD1Fr9l0DAxYrcgs
x3x67rKlN1bw5J5XLIfESO5bpRytEHyuOqvTymFMm6gHM7Tv0r7kc4kdD/kC+IWxK5aq7syhGmeR
jyMYpBIfW2uI64pq5E3sESYGrd/QJN5qTdzMUprq2S6IYrgP3xBigGwaU+pUiWnvt1Z3hEXlO/Xw
iC0YqGV35ibuvEvHI3Q8bSWl40FKts2phFzo4PDLb1D6N/Q0uWN8lP0WMFBa3tZVDHUOGGHuHJlN
94LGqR4QBGfKxpvjXFq5xlZonY5ZUWHtT4LPiHDaxMrbBJVIlRPbp0PY/5+AMfzdTfKWDDMjhU+O
kpEWyW9uPfQ5Zsr8QNJqHuvTUTiGvUM2ahqOqdGasrvpodfWty6vjyBIASfUPRdDgp7tzCxPK5si
rXBPfVGQemZhb2IF/ySHv+EwCHUsu/ESJk/qy12uedaESr4WndfKAUSWCIocCoP6/e8reje0wp/Z
w5XHvEbw8anSyu/nIyRWMKiY5QicqOkMOLZkAAumIBhVA3KaO0UOsDMO86dj8ANFr5+IQgNWmx2M
kOXLxbPW3NgpaAWHA33dx7yaQjZtcimKos399cHuVr1u6MuA7jjWZz1AJ7cG0VHxkblvVSO49+zW
L+jOh9ptJtbzIErvkwoWr/1+f83/ITxobuWiO/0IpPn8TPHi9Cc5/lnhV4elPrrn6U5iGeWzmMnt
g/633wPKWFPQWdTKtDyKCpdTpmt1Gaj5Wli0gVetGjHz9Cieafj220AWH5O6lStUart1vAGUMg7R
ORz0s1kJzxGbSHckPMiiktdwJGkz7TdA3D5wAEZGdFRlKzVFBl3Ogg3onyyrA5KWJ/jbV9wIL9Ge
AdsWjV3OgrslNfxx9H+PxWeSLrP/pWbkYUp675WfalQ9JPAyKydIwgI/QCqGa9AwkxqSx0tXDeAS
B0LXEG5weWNAjzHiMhSXqiIokls/FTtcwrP7J5cP9Ok5FTRCHAHEad2UHpX7ioUEd6EfWyTHXnzN
/lIzOcsF0hwzzlt9D2KQlasGhGOJ0Wc3mPPN4Ih+TMF2kfJzgdsP8M58f1kPa35Q52lQcfQ8McVS
ceN8xK7wosehfKEszBPYhTPNiI+LpwfAQVS2Ye13Pvj/BE11lZaIrPvYzTyURruAQyO1vyrnkN/s
Pkqj0KiUQynOXlf/Q4dyjiiaHS4XLUYlbt4EntaXRN9oYULaE3B6JnjacaL6qOMEcWLUUC9PTWCY
Lw3Yq4PIjZZgFZo6NBdUtaVYmX7mOu1IZS142NXi3HeqTdHcxaid0xa+y/hu26dD/vqFNFHg+f9M
B0MlbN8dmTlM2WkjsNY0N4Zta8MI8vYJJankR612tLCWaxyVzAaBaC5eYcxz9S87gyjvfQuzXN+S
HZou0Xy6JVrxUM2mkCSnXH1CbR4hVvz3CfzXgFGfzlhwingH5KPX+FFIGGwGbA8ylcQ8W1SFDYm4
aeHdnAGKrPvsjpqyMWRoJyVR0luW77+DQxv5zenpNjQ00OtUOttG5qmF61Fnv0K2GVW2MPZwUz9F
f/JRMu2JzASusV3f/32wyHuCpcdtrsqvf9rmgVxDK7bidsN3/TI209bCNJdMX3Y65zgi292oSmJm
+dT9zulfYd84vZiX+mim+teDvHAGxIy4b0BcfEponm3bc4tpiaXUIlfC6J5gDHEz6pZ/dCOSk0Nr
WIk/8nlsNoPZIwk/w7AOK8Ds3uScPe9Cb1yywRG2tJKDPjYoR5ho8/1a/RWfA796kbOv946bKcVa
bHwl3grhklBssvqU4nv0rugzczYklU/zNRvTTYYr1KK813PREYGkKakcOMys0sewCrcVuqkvN4ve
iH7cNLj9f5NHgoQw6oiopZAh/RSzr1x21uUSU8Xfjh57oGq1KfL9LPO6YEC94NaFT/uWFM6HGhT9
yk52KogvpsWvp6X773mzIBWP25Y96JcShdnfun2ozLGfYWg7x2Bqcrld3rKRsCyiWKAVF5Es/KfZ
v1NBSQTvAp7Zn+AX26YVBroEzBrFpf6/H898muAGTUprP1xvHTv2xvC/XI576ZKMcVanvWBD+Z3m
IfWqsh3GBoqdIB0s74Dpibt1IWZR8KoZNKpAfVFDC75c+8Blt0XXRQBl26SgSilywGWXEzFksFbP
5rkbGyyOPiorhHqG3ncsa+/d1hHw1BuxNfB9b8RTn8E28iP2mx5Q5bD/3PxqMUA1WD6Fd0WOlxfu
6rvGHSRlykHTOrznCmw+yOCdHeQRfB3APw1VsT5N1/6+fTEtMWJtfjiMvDzGhLDEspOT2CUq5MWq
4fhjJmy3gSv8PhgbpaOQPYW4hbm2DDOhVgBcAezNT+8/gkwkmPkbymRIrlE1C5m9rhJBVljqmomW
7v5dythxT2xR4KIIiYhpdQQ0wWJyPqAZmH7r+m5RvdtQe6h4LsSXvkNLHo3F+w61XoYSBFLnQGbx
3yP+5b/j5FuhYR/YYk78e7B95RksI1Q8PLrQJO75MavwctcIe7gQLbIS9vrrDkCHF2dWEmjPK9Sl
m+ICHFeC4Kqauu6tFb7pbcO0M8DT7p8o4e0lvuNKdQBNa/YM+bVpAqelpQXcdKKQkXBB6nOVU7Cc
8OhdUIwlBkXg95yqddIsa69vX1ahOsueEl4L8NhqQBV59s6luqVkHDsMtxi+XSlWM7D4koCdBhIf
aR0lzOAdv1RL3sw2Hw8dWclOi4DPE3iDyNBB/w1ljyeshelS5tComOojpfEDVMB28ftCzHa82HhX
8TPIG5wd1sEpiUKfuF+XHy0qmmyIommlRQ3c3gdjWf4zSMmSETeGEn8Wghn8toHqqexw8JT3Ipb1
9cbtLyxow076cBQooYGVL+MWikf3Rv2fpUkTsVdJRVAAyvgRxQXTz/tLF8CIS2GI2ucvZFTrVv92
t/qoH28FzoAVTI+TrVz7SlVUqUwiDtiSw3zF41ucs9ERSzBZAujmFzrkGAnKAp32Z4laeHm6S/gz
+sd+8H5B7JeUuN05L+aLK0f18m2k32x9clgylfVpKASZXYhNwLwzwwu+w8P1pJeWuwvtRflS939R
4b/B3MGFG6zXIQpeYZeKeSxeSjF0a9Z7aQB064sAGDiJfmTMB2G6Y10rVFQuOFmSLTC87uq388T+
jQkg1/L5lWeR/9xSkMJejV0Y4NLAnWaj5mnPub0fQXMQLLWpgqe+o1hDDSg2zN1/ge+3Zu7R10tB
ZeawNgYIFMPuRKG7FxqGdlaib9f1ayadGw+rd65lloeTNeh6zMztSZhoLgXc7RvCxCcV24puvfYw
Of9+oqd0++CYf6K/9Lr7pJe/8wEe0kUGk8OwCv2wzi6i4B92mvoGlLH3q5EOS6SzPfDvAj0h6xV1
ciX5KTBZRK/YqJRK7G7pYAlepGafGsfXLHroPNEVlcNplyirNufbpb/oF+U0dMRWgJyHeUME8bnd
zDPvcO6ZtCg9oWmMtcr3UvZhUIil5GSDC/E5SQIFijaxAj0+0mBLZzE62vY0iZhKfNi5MRkf8gKP
TVRjntogCtwARD76xRqLkSzOqJY1Cwcm9r1H2bb/KXeE8sRlyAhA5d6lZZOKzWuPIXkZ7wJuSO1s
n8h6k6Ff0DwG3g2U3/0BvrJiMsw3TQBRkOEjMj3KAZlkZCCsLLldV0Krvoc9P2/Bh9/IKWmLAvj+
Tk3tisJnN7V3ckBgAlYe5cWVwzlMYaTuYoqr6pZa4KNUSMXnWARnoLJuUowMzwTrvEJyJAVBsrG6
MSK1/pHw5/KX834XdXYCS97iSp/G+iJjkStARr/WDLUlZWPnWSJ9mAs2vVj0L59ZAuQOdVEwZWMN
OqT3xXsxIKih5r6ny6adNyz99ZZCABmwtBBHfq4PV4f4QDUUaDAc6rEB0CWHQvQ/9yG8j3H4Ho31
28y1HiWQ3zSAhZXJlwEU6nM1UqhyHepNk0HeqT3n0Yj4H0Bkxc/UEvibsOOJ335vrM1ePMUAUidj
Fxwrzu8xUQptefr+SRJsXCYQCmX2Y/KFtK49g3ejOt8ipOq/bFBf40vBqujh6Oj320o/JlpRyIRF
L+GkZ5Y2m+2MyteOI93DNoTLBfApY8KDL6ikiJ/6qwy39D+l5NlMkMoz2M1gAY9BNYuqKW7CqS9H
qzwzbcDrgOd15RCsmiLpbn1JsCSX/4fYTaz45nwhClK2Kt4xdti0gWoo5tBSP/FtQmJfDGg59OOr
6f7jMCHSLV8pp3uu6TvlgdTl4Vht66Z2hrpOjOSwrUQ5ngCRhBs7Uqc72fL7C5xybODypM5xBfbG
y1lcwywhFV8FBx4KhEVF2a5c+Kc1VdSG/df37768xByvOb8DoiTzKy8ZGAOOx7ifHM0nmuY8SgYK
0LTxsA8/6b7LCWS0KHNmAdb3N2f0RLZQEiEzx8Xp6KuzpHiAQToewWKOmPp0IqvpnxHzUL1bElVE
Y0VYBltI/yrfJdTBDY54pLUZbKCPLl6OlMDjFGucB5YSkJhwdc2cp5qLxNU7F6pGL6Q6v3zy7VHy
Q0DbD/yEGz6kWe4SLQ2eaV1Yn/9L7MIFPyIz9KBL0NXPsucjgfCGrMpNBLYYL5aMlQGYlaof6G0V
95e4HASA0vT/iq2SYpcZIrB1FBQRPACGeyqW2mgm2cBZOL8WK9hJzrP/H6JodF4UyDDMDuhHkRrq
86qtw/P5HuHqV0l7qe48viB43oZly1bQNzilv3px9mt5+t9ETSURB0ihoeCGOdm1sqffI+b+PFLQ
3ZzgCwbPKoh/cOfswUfcAcEt0er3JXzfssTyPlSWfTjjrOhDf4Bh9TaDkg+08CWcaILdA/WFoJo6
YSwMuG3A4mx6uV4MyQ7GKWEJpHDRZsxRWpf4jXGkro7NUwvf4Z5s1k/SludifKhK2dJNe1YAexYk
gSsegDx2zEuVcu6vo7/k+LMbFjWTLgwifrDLFnC6BpqJLSExgBLwtS44MRwieK9LCBnjMA7JXZKN
tIIeEzwsvqJKvl7qLpgenda0PUlYZe76dMo8Bp8lFHqoHpJ3qsARZi+KolKQQBFpmL0a0Xn4zQon
RRhXtHLgcr0dViI7BjAwnVkuSimnFkESAT+KR5f1oe3ZHb2Fqelx0b2Q9T8FNw6SJ5elBoG5xy5G
MySEzOrZ1sXz87s7wfRLkay/ySJ5Kvm7HccXq4QyoDD+mcPGVkqfEiltMWo1gfu6slYeEe0xoD6s
vutMpgZCiugUKps8MUamGl29JC594LzO9Le9+4xgCAFsG5O/kumUoFaZ0GjbHUIratmtVDZ6BtyZ
rLKI3ug1wf1ktukQb5VhFRy0F4a/OAEzXqxaERKj6l/5xcnsTCr5RwXkYOrCrxyPeGgZfM+2Jpd4
7prFQ1eL08r1BCD+PaohZdgjVKi/sIk0NnUGBCZKorMeRvSXki8Qjd0BSJEBzYxawy3r1Tvi5Zjc
YoCmoXZNyjq5pFvuKzEkKvFLPwadIlO8NXgLK3B+OiaA7LlBd8iOkWowQkqbrbImwx7hckCdJL+t
yElLAY9qUSYCdhP4YDRJTMvh3/PjwCUGY/fyc8/I89T9vULqg9vfrkeaWtGTEbkNsJq9nCmmd65j
T4bhYCkoVNpsii4Y5qLYETEALu1wO+UdXbOQy7GtggABne7acU7OAYlAF9LUwPFYahK/yRjVNgDM
9sQuN36zeqfSzDQf9hbV7c5N7ZbFN8CSwkj78Qv8fE1EUYo5C++o83KF4Qq/m/ouVfkoWYKEclXP
cC4ttYFs1F7NGKbD90hnDvE0tTc7A7JtQ+i5Ok2K4q33GX22nuMPvFxOegP7DIXN1lH3aw+qfmOZ
iV6egTGN1uQKuijVwq1WL0pUk+Sn81getfuxzVBNzrSOu/dl+1kzmb+YOSeXelB8518U8AWrfVaa
3Ic4T4Y+VaoVlqtRFL2wIGJg9up0xeBrzI89QdmXJ51Eqmd4gKjr/JtUf+qXPpzzStRh0L3bL7EJ
3MT5kQ5f32PXxWkEyFVM/KkTxPY51T7ElCceJ/yspDSfLeI6TnxTfxRSKPMwphIYUB8XEC98ovW9
kw3lmZ1/CRD8pIW5NxSiuvk1bbDIaO/zTPgJX3xyRMBYF8r4rHq7MXXFkbG2b5fTI1Be5w+d8nOz
XtrPWIT03Jd5VS3hqbdbe5Ykyok0TV2QdytfJ0iS6gG5nD7EG9U5oZq9wrjpN0zwr4q4ReAuop5A
KTYWp5cKTaT3MSmCboUE88c8Q95g6H3j1/qCbEI++BYvu/Gf+8NAe9hmo7YKdFmDdAxBlojXzIEX
zypQ0raDMYZL6p7OADE7rO2sDod5Yqry0sAjHcohozSmh6t06aol+7aPpmlQoeEBVtKC7lKaz8Sy
oOyAb8cRPh4P3/QCtVAENRIYnwwI2YPqlhstJVu6N41wrtjomZP1oHz9hIgs9LnJaXi9D1GdT8Lk
tBbFXXq1YxZAJQv3ORd0iKMZdBNj2znqAj9HQo1+37biYb7szeuEJwT9zA0CzWnqOb26xyaRDauN
NW96yIi2ksNkBbFFmO9yWULOW8wm8Gwz39wmdJtikIdIrET8QfnB8Xt8N/j6BkwYha/3T9S9EEy4
dZ9S+qoOUZCkiusGrt/mvYu2q4887cAkDsOVN4tA/4iZt/jgs5yx5M78N022u2Wy7yNL7RNMx6SM
hGgcBQyqdBRqth5BrTC8D7NZ0pjHSA16rdo1eevKn0+JsQa4y1g9JOL4mmAJ0+p+rLGbz/wrj7af
QijhPxkWjIW6BkJ07LEVCVAbn/0iUCzWUxV3B9I267tMwRHjZ5cY9+SxJMOLjceFEQ6yOsHGIe+G
5x9tZqDIwAEZvkOtkVXeGFythKzhDkJmR5neteRKYBmyxzJYoODFlywyI/7O4QN2Vf5LcpDH5223
APlXqouoIRrKT/nhx2CPo46N5ysbo7lkr9JWzpG4PJG9Sbo8lLvIK65pmaqjg5CsBL1hjiEwueqE
Jam1JiaCQtVw4nB7A1guINufHpU7h6ZP6mvqpjvxidlDJe8HfCcm9H9lZeZfF1i55kOswOd2e8Or
VLjIL1+V7xkfp2AuKdRhJSsKssQ+9Gd2edhTjDmx9mmreJ2nbJ0+A2xY22OJUJrNKQPTdSX19TAU
s5Fu/7VU/nSVZ6hUxK8KRw0YHXR/HPe2odayhKVTSwR5NMy/BwxjIVrr9fpU2uU9QbciZ17CDuOj
ALbkGAtg7qXCTOlEpwAp4+N11im1OwRnogngdnzMoiHupR9En1MLzUx5ZSGR7d6DcMp7y5If3GRT
f0hopKp9nn9Nz/cPA0RaPDeKVQux4xykguMsiJoegNRdMZRpN7159oTt4d0WGXPsiY4hYfeKv9cn
wXxrfyYEeBoKVdYbWhoxhjVx7G06XEYO1HnBQgfIzDuQAI2SAzMjlZF8jpvGkzPwRcOtV4lp6ThS
yjEWvR28eaU6+IHMH5HS6LPlIEL1rMN9vxNsP3uKOOebTU6oNSmHlZL0m6aKYylx56g1tmbE/0+d
ejZplNBq/teTwJcACvKfKdFMVvgiMtq6m2RNmoK0mTjryPTLEJPs5gC2R6HSYTvVrtsZUiKC+lAY
ZGSX91DVdMMRHIbZvsywY+nLaoCIsjT7od7+73t2MHo5OIvvzLw63uTeD+U6fmkfXsA5KouAy9HE
ff78XUahbwCSj4nc+j+WTRnOCgj1mGmBkjopK5GR6p/v9j/v/SUywElZYAcawgJHlBEs4z3r+Dz1
6GU4So9/SSzVQL7Dj9ZXhiv4nQBfAmj1vy/s26OK0jBiMklk9tHRkrAxuL9DXxH2fOLgEgbsiJDf
tAX4ddXdpuW+wuZERSYCBVPyMG+kffgY+Dhd5id2ICO+gEpNg60fuy4E4u6fvfJwJI3psgw68VXi
H6UY4dkTHMvc8JVGWsGHlNbXWf2X9mMOR8eROWp30rmET6oXnVbZYzdTTCLg4B0UYfJ4QuzemkSo
pOT/PWiE6ojsCTot2GQCvsetc9NSFgN2SZWH69iKenWszxNzwx0kpcbR91QXF6SWL0PCR58/qdWv
WOp+fDmg24nEOrqNd6rWGxNsOzdA5ppgRRmRd3ihekpYIJwjyhcmbEC6QGyVhfPDjMo9DnehdBp3
EGgwCuGNxsumnIZOZRbPy467P16PRyGTRjyCdqkU8KrSABmbdZXtsfumHNaRyxL2vLMZ5ntbWG3d
iRoKzuhBqYLFPO0UL1RZHQIzkS0WlxMShbbIG1GD7Z2ioH7GgWdKCfsFXm+Dd5ghWUEQi7CSQqwg
lw/mQt3PbR1Si3ww0xD3gV5US7aYQr8yDDTuHGjlp3bjjhFtWoTtWApjye34IoxoTYEudRyjwDfx
Cj6IcXIFkchStZrLm27NGJM4Yy2MB1rfGZcjqA0K0f/joJUsaphO9AcikCSfxGs6bucf4knKycSB
HHVa6fFmZRDELbZCwW02b6oSubj226JdIeLAlN2iToAyXsMZTeL9zb5okFUlp55f3HVNtSVtoIWy
dBFm1adnQ3FcCpbpx/e7uDFZzK906sCw+qxAixQ/Pwesmd2cHwE2+N3JndMb4FiZDWm+IKNlVwR7
0nZF3SHc6ySlCHosrt9Rsn9b1XOMK6wXhjHh22GPNcSWWYoN61Ix1WrvRUbX3XyVaiyQsjVMV2uy
MgUMebrgtBVs4T8g1fwzOkzN+o/WUo744z+0gLEnSJWedcDmI0TSWK2ID6lPNw0XNZ7ZgJ6Sd9U3
aJFn8R9ocOSTA/ljvgLVO+Km1H3EQcUH0sAR5AZacu4Ui9se5Klpu/cOWmDqF1Q75Hy8O6mXBNTA
6q9UYrLW7XPDWml6GFO5JId6VbFYnbvywg2fhh1Ggliq7vQvqr0ihdEDc4YcmrNB4X7sKEEHMKHt
7BTYBI0yG+ZuvFdt1YcS8qppzJ3K25qrJbmV/iNVepUHU/i7ZxlKcTQimRnu7Iv+R3k4D4/MPRaJ
cJiZApHCIqwyI9SJOStmIsKyR1t93JkjxhEWB4umnrje5DXzTg3tzWxqajCF67KmkkkyZMwan076
fruZlNajegU8+HUmoZTE9WF3RALB8Br4llhwnFeo2nE7gCVUz5MfhyIIcy8qj6CLzUWgTC933pEJ
MXSKS3nvgLkl1R9MDSOX8JHCPWCHqKAiajazd6aAXzXsBsau95zAcmwTNk0Jonai548aRn7+M6rL
2c1wVWbEm2rqN/mngTyHMciOb29h6XvJU/2q/bEeGVT6GzfEq0gL77kb1xilwAp1RwsN0Apz2GlW
V9wx7Z/ZJIhCRGO5ZlBSBwIltMyE/L9EIn0y9U/n3g5y+8mbStXCKak+2jDnpzLVppgm8eBmpTno
1UwB1gBtd/gC5cNGBIWX54slKjmz90mOpNhz8xIWHQggrR/AlHQONS+q6qrG8ojLpv2E4cpNRLfi
Ru+uiOHRtiXpqiQ+zPhketT2ddxfrznNLmaWwpenFj72jqW2Ec5LSy0IEzP7cr5RcYGfE6T2CpZu
ExRrNwkLVKbCoBIGXJebkpDYhMidifjM0uvp42Ytqav0TI71SDz5/1G2JCHJFbhVLpDMpvBRZ5tg
HjdoQCRM74OwpW4SuQfJdedSVRHeh//7U219/S/zwI3PDkM+qEjZzCe5ntaZeltclwZcE5C506Ee
7ApXEjH1sD28EqseufZo6nD0P9rA9dOEkbY00A75Tdu0ju79cO5rf2CspOirBgpCEg9t7CCIDXDq
Z3OYmh4XiZwX4To4Gc5zopQFURi8kVGSml+uPTj5vvAeB60nnFI6jY6kI07gEmjSvswQ+cqXYbPL
wdaE+7n+Wd/38D2soK89ruMH48vGmqbQ7oviWMT7NFNpWDzzWVGqHnAdLg8AvneJN7FhDhpbnznD
jD1Uu2H7xjtA9qpTVAGVmyINEJynG7fmPO8Ha9BPdTONO4jMiknsO10ZDB9kxmf030217QBVXkMG
70mBwyDvIb0f+TDnkGiLiPkMbNNa9L4GzkCO5n8xN0BzSs4Ri91+jkiKdPaH1aj/Iew6S3m0Bkoj
gdkRkRuwyV6wx1OZ8tLw+P8T1CZLgP5Owwj5lTVcdumeF31VQesyIR5koU2R8erwG83aQxmE7QyC
LhfFETEiGydPM7lgHwnhKNhK4/3oyJJuXRTKESl39dgU1ajH86vHZSaSgNGf2/fCbyoPN5LoaX15
KMjfXpe3lWh/1ckRDjT0P741xxuuTMdZHFqGjX7tECfGO3YjTnYJjuuAS9z8PlWOXgoXlZAKsxyc
+fKrAVJ1tsuvQJ9/JhZP2qwldLVKLq+6DWWne30qrmbHhdFSc+8ZNHc7U+P9K4sQ12+hfIura4BQ
VOoxyAMcezSkykDp351HamrhsMQ7H2Mww1CWQ0S6KQUQvEO2KvaA9UtQdmW85HGs4DMKYhGPwnv2
IekINeAczvUcgbQ7wyEoY2He9+pSf3jXEoR0pPf7RzsLTwPBheQOKMia2Vcwr47QJHwB2jS9GsHL
dCK2P3ebIpsC+Jr+fm4l5CpGp8JO6trgZ+zQuaYgPL1KXdECgD3uENvQp1R0P0O0wQkQN1Fd+A50
oRZLgDh+csT5xVfnAUL3EfIQLCsfA5OJRk01fXPJllUjbgnCIi9z0wpQNQcSwN0o0k6R6fMCa8tN
5AsV/Up6g+1wK0wUJ9sptp4r4LF58rsjQ9fZfn5RBcZbObNLY1GgnsQIwcXOfNZi9Y34jr07NarH
c557VgI6USCkoMs/ve6Wj2vPKWnjnKoYuQAt0XSbPt+7cR8bH8ahmPgeN6ME0MlFwIpnYGCV1rBO
xZcWd2oKIhcn9udOTnViQ3BDJMsvvqBuF/w5lTPrAiihoUvCX6+PJDSJWIDv2gsGILKz1Vt1HBxG
1bM6Jy5GmMMknTttZuoBzqal/39+mADOG41b5gph133nNlp1jylHpXsYMbOw8I9f9nOxnDc2rDVt
dAi+GgGYf0fOGHvfmeuR/dl8g3LnYiaydGxiDUWWV4hZe72CAB7GpsTPOS45zhIXkF8IOZ2wFOWC
/01eGCFM59BZ4A7qRwU8oIWvRzRQZXZ748lqWWa7X7e0AgmkDzq38+ctE/fXojkzq7zSsBgU8zdx
ZHiufIJsh/55yiLwlS3FHpqr2Rv9kqDbh36HB8S/XBWcfMh7oHp2beU4LM14dTmMscs9QSTXd0c/
D2RutFItMDZY9O5/g5yr5jNUoS5ncsShdMVVEu9W3IKbFh2fW8EAzCY4JszsuA4UflXSzHQn/xiB
uxv3CF3M8H2vGz8SH4sXKmCU6erwQihB9rtYtkzjnkkuPxSlRAT9foLwjNjN6SfnF+Bhk8s3yKmh
oSIerKn55VCuyXxoEgw4dM8Nj8pbf8n9CyWTSJbEaq/FO/Rr8xY/QlsKZe5OcBAX4X0C+6VgZdlX
9MJUD+3JGS55tG+oi5EaTqR0qg/VpA5bCn1gdnDF2rk9nJf3Uo3k1baqtZFtBXxcuqd9tAQ150pX
krN9pQfeVvAuiSaWP4eXYxDRK5o5SHVf1nfHpsbCNx2XAr401AqM377TJ83nXE1jO3K5DiGQuKi4
/F/5giRfc8U0PSmGrxaWDKganS+BO0QqZZzxEn3nFMqhJ5Nd8NFJu0er5FSC5KvvI10rY+akNt1s
VxQbBvwXOtK+JDWa9CNYZJg5Mb/a3sv4Me1aQ2sO/KDHa+QfwKZ0MsW4iOtSddefAhmZ6OlRwEkg
svtNOhsFHy1Byu6EIxYrrlyTANMvFXlltyRIiAtgyvftZ9urEC7pn9U2FlfqGGvfeKHWa0d84NYm
qD8TQm3dKHsF4/1ZgkkA0o2MkUBE6xCf7xBSoeg3wlXi0APgwBwfxXmmPtVsXj46QtkFkNHlOZ00
scuvdb3/JdaSWx+yFIo72GHO533Wp12fkYIQWp5LF7kzJxhugcalbeI0kmuHfvFfHDEEUzWTVJhh
lkTA3tpqhuTR62DvXvgoSCX4bhNB/nVYz7ZtdtJTCgA9y5TG/D/e23sj9UApmpJ8XCnbWyWVOBl+
SW8DdCozkdmg02ySdO6SSUUyDbnkd+2kUJcT7TzR8rnO0xKPGcsZHZXcsXq2LG5fEAe9cK358suR
zGY3C2PiSsEq2Luk95FSNfTn2CX8CmfmndOfu7LTUbqy1z++4wV6PsDMky3TDhfLJcGvxQ6PfzT1
bfeGGAHBauTqGLJJ712S0e76WBdtEMv9FqAzzSi8GuPF4cPXA5R+Y//naq4GBGP9zJM8PydTTbcp
+rnpCsd6kmUDONdiR2242HJj4SksLPXE0vBlDYS/rvo1Bu7s9u1prmUzi78Lj/V3ZBLnN1AvJ8NG
3PwglQN2HpUWJGZmh99BEc/pXzDTCuSebrh1Akq/1n+BREei3sScmMWZuRVPgilOMrmFF7iGQzzZ
WDQvfC/v85Gfe8y5aiIzHLFdc5W2JvZbURdBzDjdjqh1rBLdT9PGXYMMoVaply+A1umHPlpl75p+
fA7TXYZExCj0UBHIRag7McICl+wTIWjU8KoBoom0/VKU+fzGKzd7fCpdW8Q/OfzYtuwSBiAzCy1Y
nzssOApahGMMdaXfPo9wehaD6zGIOX7yKpe6hZnZat0X5UsoatezE9xjlCLWCjJe/x77zLdJWbRK
rmiNOwPier0jAeE/ZJtjN5X+7dyqsReJB/hQRpx4A/Z4sMFCuvcsj+wTmiw0kZBf51P41wNJC9re
UDkb579Iv6eTBldWWMSt8tiwHAa8FTMCpCOI9HU87vqbImPnFehjPHXWvRUvoZvuSb/cF/C3oQ+j
yyDkE+CHwvA9Wesg0Cwib3GsAlaU5fCH1Mp0LJof7oOArHMNpGQ5kUMPzqGWAe2xbyWZ50uPJS0T
MXkBXZU5IHVH/maUMfw0o5F3tcc0xq15wI6GjRWmpKLcyvrt/4oNbR3roOzcazQeN147FF15ys2b
OnltBYk41VCSluNxF4flRcFHSjkGgdVEAW5koypUPZbSI+jRztIHrgLin3toduHiTKPDd+0xNx5X
+zr/wA5OQ6U3QEoKYH8UUWwYyGG39xgeBZa+Xi+EN7Qyy/E/mdLHEqVo3MGyHTw/jyUL073GAtvc
eGyEoRlU/BUiRdhI0AU7tyWosf527WRtJk4ia0AcPws0oIOy+jVtohhQH0lb5PKe0j3OYCl43+dU
2T9PF8lcnPYU0etO8MqGw6YhuTOqe28yiivnE3gQtBqZjejAf7VM4nxl/EkZdGTktb8wvcG3XrtI
TTmJyF89JlUwcQRgcfruTx/ORhW/WthWr6wPofMkqRP3ZmN83kJJ/jP2NjWuZSYZJ96JQ9Gh48bk
hpY8Q07gvt1Pab6PS+nbUXIkNB4ikyGcSF0Yhyhi5Vj8tubXXdIprAA95gW9nv580EsHpGfY+TxX
S3YAwXaA7UKPp8vI4Mxuvg2dKyQ0bWBM0OOZgNEgWiW2ulBZKHZXInXrKS8kmEBzIlzaTMyNSfZ2
Y0GhqX1hTCZcsx8ZMG7JChc4UFwz1pZrQi6AMmNfLBhT+MXJWrr4+Q4aEySQy144r5mGAo22aAb6
Cel+19D4pDJSe/A1YsL55doOQ9E/JoXzNHBYY31nvw6Bld2QM1e+y281T2rcYsaLA8uBe6+KELOV
wTGIyDFdCFtu8YWsUkvHO0gpp6y2XuAcidlIO1oE1fgvkSRkIqaR9h/ccZmqu/hbSxm7Fck+r9gt
cic0eY/qdAbi1sWudT5sS7+k6oNkjjljGtIk2btSfNxn6Whk66oCLcelhSlWQ64uO/OX5AQhaxLk
DM2REAceVtJryaHPNrJ8nNQD5DqQIp9lbY/B+Sa1FSIrplTq4LtYiF9qwGSDqX1yizp3tdbJkAFG
wuPuXnqkHOiQ97sORxtgKX+qUjOBDMKNxi5fCST/bZiS6ErSdtsw+O8V6lgi3DYMKlYFpSzICrS+
J3Cooxa0x0i0c/Euqs2s6yLmphgSFBNG8cMzTeuR9j2USxMSRD7NMeW0K8axqAMflujDnVdYTjfa
en0M+Zqo8yCaysXTzrEm7jyHTCHI4PhYeoocHUpMrj8PaWj3TCb3o0CdrT4g6PRZR6Cl41lmX6Kk
L3OHll9PRTfxs1AcoQtvtZQMyQ/pS1yJ/D2KDPpkDBIvp6ffrJQeikPll5XDLiBAsZHOUojHz15Q
VlMx5K00pWkjIs+ms3CewUSwnrTG9RlzG37GLAINOD4AzOj1q4fvoPlsZ4z3gMZu0LNf6oaARBB6
4MSu4LaB4+JQhgkiV6MAb/nYK6kvdaL7m6Cqn+iGTfjFT2RDAO9B8PQ1e4mgZerr2DfQPYylZ9hP
bLU3MF10nmpFnJJH712sSTLe1r/Z+skJB6LbHLzEZ4LLHtUYdGSkXz81O7uGcaaj5IWBP5YBQsN8
bqa/CuI5yP9xXKi3o0BjVuZERm3frVUffBRCOr/2rD4e5QCfUGAlHDg/RY1CZ/V9HXDJQIlXrsZs
onJnDAsK490Y6Pv+qoOb1Fqy3WNq0v0cZUUiITp+Ox/MjsKmQYDzK31GCN3EMWRDWs/9ybCeRuHk
ybADfeKDSlzFZJnXwsDbtKpHHVNypg9xOizDDhc4FK17WQMMdKqc9DyPXx7o2hX+dfmX2LLGvDmU
s+YU2jtOAxKkwB92hQlr+RfKRi1sMOobqaUpTjlg0aw9BFNqYD8p3TCavm25O0V6NYLvDhGddF42
Pdza6edgEaz+4UjVcxco82QbXWsVBFFuJXJ5fXPKsQstQzyFUGXZAoSGuld8uoiJ7EyjAZHiuhcI
e8/nrXuIGq0mAJb7A5sPy87Ga5O+NHijgJg+zqSUbkF/J8xBtSNuBZ2jLl6RgQDG/tpnj/7nNMDi
8lE5dQK1dgHHFfCkOCa2Q3rCJz+Qk/AGDNcNamlmeHrnr7Vy6nC+tKIiU/nZdxnlsjPSFbMPG5Vo
Ty5c71PYteP0NZLoL0LpGAFjbbPevHKmKHnQU4Xzf36+WnK8HpfziTmv4iOWaOzzcx9LOWrIFihR
8HlA+/P9b6NNtgA0I+k/zdD5ThLpwg3kvJUldzGsDL106m8D/jPJTKsV2v9xd7MNUTEh2ZBten5e
U0/LB2bhTBoxJaEwaIPWm3dypK7HCjqTWvAvPG2cUM4q2dbXVfoFaQM3XSlioyLFyl4bKKzq6zFu
eppio6GQlRdRvs0ECI7lppryelNAbUJkiUiyt5PXiwxOLgr3NOaMAk1DdRzCxpU3Cioym9oEKRAt
n6a7kaXsq0kaQFQIYj/juPCiYj81pcaL21CQ1uNR22j2HVQEaqCbBkNrlNGpp11DmXdkriefgJPY
nmtbAnml3nGsIsL2RxLpTaA2y3NuRYfkTY5pcR4FkoJbnGyFuMeC+2ZKq6qT5BbbkyuOThRz6SiP
1R03LPzoGP+HKw/0pPn6h7D0fPXBNeDsu0sc5DT2Mx7cIp1tzgV1GXESgF4f8grruJyp/idZ+cns
XhSFy+1Nb9MzYHjANuK3vsqy39DjKYUq4qCEfCSethkqoQ197TBOusOEXngICaPwNar2Tz+RGN/F
Lb2N4c292j/A6RwI0ZMQj7SXmvgcXJ05+etCNJyjlxGt+YVvUVzDIry1oP2sWHrbXw6l5mmVEl67
fhk/z5nZlcdyupQC4+B0ylkllXW9k4RIygbgDPowQjKOUiQ8m/vL2ZqHVaFgDceg4knxCdtCkgUr
rIJdX8GKXOl7SRZb0FmrYUE13SUm+rXGYF4Cf87y2LuirlACXfZUwyeyVLiyY7AbsCOPndjpxqwk
nxqzoy6VjIZcz4zKdt5qwJ4sPz3AsemeVSaw7OIoxC7oB+JWXDfgfC7JqsBs5SGR+n3TzfJ8ltdy
tRF65Cf9DGSHKFT2bpo3tCtEv6tkxzWsbxf/nZHFBILSIf8ytvcu+GVB72+g5YNMrN2BTYM2DrsB
XQTK0OOhPq0sTXJ+pdSP2f6ApSxCQNGbC4M7QFVkev8HDSIVMe+eQV0K8M4lMzog+7RGCqoGlbvm
hNS/LtzC2lGKT7DytHMuSTk3tCHt83C7aHJ6IxnoNifw7Ho+XdtrzVhD6yDGbks6X4Nbfm6YoQcG
vAD5zIh35W4qIIHSn5wFTbjHAOWZVXPcG4gmIiHKlkOvzagE6SzuXjPD9PXM9uahF16KRNiemyyw
sSvTZYHAV6rHmiCYuRgPbuODwDevIrHb/MApnV/qgCsm5blMn2/Xb5KGQkSZzIMI2Fd5+/1tVnAg
ebi6NONxKQoAUX5MlJgI+0joznRYgXKUbhc12xWUn6+PD/roSR1+W3CJYFWWcNi8kq4AqY+oonfw
aVCvtRlrFZWG2J3+vdNCQGDgFSQFyY9aQCWvBaWtRd9IFan31CSKnn5H/TS6GZhZ7bSV83bz32fz
4ID6y2Tas/PYDG4Xl01byd3vmu+YyuNCN6qpn57hXv+uiaKFDv8Wfurhr7UDuVo5Z0PD9M0uw/i/
0Q14TT0HdvGggUvyXvmRMKr7o+BHjvhkWStCRTscAi17rcAOB2/cqIpEMMjbv+lpV4qAWvs+BbLt
+rVIkB+FBjUnJXhIxB7MOc0ANRci7uxRbD/Wl9srGmM57rCogbVCc6P/TlOBxf/ZHwyagCLkqyu1
hgL/BOcNVcc6omKmcBg+8e+s5l9hMJmbQhsbvvGKpv+ym8rmmaXpBcsJvRdpBz73+49MjKJNwPYP
DkcD7gR3pe+XzgtW2z95GiZQSwAcWslGgtMgONnRe1k+HKDRnfs13vZfnsrwpSPLd6IiCa96+oWj
4yI09LGSftB7dPzl+HTBplqAgqK8DTVIl1oNp9zftynBvJCBYsMgaXATZQHhOxDCDP9JdNkrDAQx
CTDbuFF2xsNrEowjYUBzOxU2u3yV29bZmk0KYn71aB2Opsv7vOKmqcDUszwqBYBL89VIlpF2n8Oh
6A6C1A1RRHtNga5aT2HnFqsL99Wf2ivphe3PB7Oqnm27znZ3/Wr9+HVk9DlnbJ5zFgMBiEgHIrM3
5Zo0C35mtyHAjDdE0PZ3/CRy4w1FWlSBDRjvioZbkKd9bXQS/NajEUji+cTDYaR9jzbK99FJaphI
Vp4o1EJfYJozLAFDUE2INl46+6B/s3aRpTY/5yZsCjSIgMdEkF9xKcyFxz/+iPUs424XvPsZYgGH
il5S8cQ/8IaFI+7+AmYhn2CxQ0bagL7vEjEWv+5DmhVxku7AyTjRFoTH0QhWqhyXCuxAn79ZVDHd
c/PQGfoi+uqLQTj5cgpSnRk+CbJVRJHO7xDLhx2F9Tyg4qldgsoHWFZwudw7Q11TesgwWuPhF++R
MWfigbj1iLlTnw3zGcqV2FLnAOAUoIZDTxdJv0vwWBK3NSIs0o8S2QA44CBLF0mI5ljqY9x4PxD3
vC7uVt2AwHANjtx4T7eEKe3kYvAQh2t0wYuCGu7al/938gfjmuTku+ySPJhx5xs7XIyB+vz5dVFg
2JefdpUkP+jlBLuN7RiDJSPRyDjTUc5myKC75OEXOoE6KLlc1BDAyYse92shicRuI6ExpznFLmlr
JfSRZAj2yAbgGn/8fEGmsOAvI3P1nPKulWy6eyy3RIWYnfoOBjVfEHkmAXtiuu9FZsprqILfO4BW
9x8zPf01bTFu++5CwtF5bpob3iA9heAUGUCxMkOCF01KWgmtnpYlDUWp1nbopZ4BvTtOC7GSXcQZ
7quM/WELhyDGRt2pXpnOLmu6u94YZqOhN+qWBYD0Hf/ZvWb4h3bPJUkV0ECmZlwhkBoyXoNOIbfV
PbsgPtjr/5icdl9mF1HP5d8kHa2K4K5HrouWJSVsXFvwmVg0eVNi8RibOTheViyPkdHaxVlfFxc1
EXvZKhOpB1Bouz2VYnPnbFFA0h4jhQC7DGCPF4yElt2YlY9DqGPN2IpGc/CCIOQsKnou75RuXzIs
HHVonp1Ajmk32wwur4xn0xxCQZEWkbquOOoEaqK0aDQ++wa7HmiMcGNHMl+onn7yPYIuXw8ZU3wB
PCWaTEEOF7So+K12lnedQPYa5aCfHXy544YEk0xlhEGqzSUDRh6BlxkF/cH5GHasX39XTie39soW
Hbjzpm/5mrqkxz7ddqheoWXeVakUbxKk1pMq51cXvf5LMoH9PTShVZeLhfKQRReBAkH+IGgfoFPm
iwyeB+QxSwyNjT8t9grAO0mAgFm3OM3K+tvONP/MN7UeSEI7uj5ECf8r2U9s+IVbWDqUv+KytoFx
yP/NUjSAEGYDPu0V1nFBHwYovAGW9SIJaTSmp0JeRnoKLVdNRlDO32Ze0XZKUor0JXp5+vKw0/vS
Q9vxCG25n6KWs5Hg1LUctEXyDpyp52SqkkLhRp/Tl5iXa3JVlJGLBGEYmwTrxswwfSR7zkfgwbHH
fqvD0lNtzahUIp8gxzImN6prao5B/zwZYTTJyQfLX8w1ax09fTN0tb2H0QRW8+GXCLAZg3K8HhYy
7ZAWytCBA3GTA9/dEbEyLvHDOmbAs4eYaK2oZtsVZs2oizRFwCd0Da/alXGpve77W9Y9CPlUB/1y
oC9zqum+GEe4fKzCVv6/YrqbbffPh50dUtUS5vevUmfJYeFJCBzIjO842HHNy/5HBnyOCRjp3szn
yahdWN1HX85PRgmtYJPw4QFLCg4pUMfj1nRpyLvlEJ4BhkHFGYbF+6iipYVaJ0FJFsYQ2Ur6COu6
vGMbzmNUhGuy6sY1xa5fUQYfMsmAMTeRc5gTKhFLPawfYgnQgnNUSu0lU2fWJ25bIhVis4BKDvnS
uAx4MiI+7HzF04Tg7ZCdDeL7tf1LSAIrFOD76jxWY7wQIYvd35EjzoYKv6DgYCQ2Lmm96s037y9v
zur8PzR9RE2aQ9r5h4vtNZKyLXgqgWMPdu2NMLkkgqKNGQJS1Gq9KnjWciF67E8qArxDySaEuSLg
eFdFXnr8lgubMKDUW7AayPTUtmRZej9Tubng8GcMB/ogx2BLcg+J0NeGyJkZbEdvb1mssamgZEO7
4rYVZGCwU+3In3cb0L4f2FGUdeSOKfFJkSeVYWrk6YAAlZMjTSr5/XaYkOmy02bM7ZnGxcTdzpbn
VyUduDUPozO98MHPE73udPK2i1LuVPoGAA3X8OVo1UHD8rToOPc+OdavAcjyFzvmlkSfb3bW1vrH
B5KJqbmV+E0BzRXLpjh2+WXidTfLHm23C7q9UeiFslmWN6n0MLbaYChONkvIcORDTh0L+D+1oYTt
N8OqaZ0umv7203Vc5qYMBHlFh4KD3L2JUb19GD/2+e5EDGegNDEQ8vf50defibgYqWoycrqIbyUV
WlnrIHGt83Emibf6bwSjNIRUi5HlbGFQtj+202jK2Zl55lfzvifZZGIyKuuXmUKsADAYtHEisV8r
ksKd3kPO1KbFLsPvILyjmaEkLWxof4ggQlEmv5hvbABeUXusgQ2CiGwQpri5P7CK8/oy9DP0BegK
DuDm6+bt9Fr4UQO/v4gRmvERvtTuyTZ3QVdoxXx3E3ox7haAcjwm+u/TM7x4eIcfw4EJFCPHfLer
fAi+r0KkgGnN+2VqqoF4wRzM5Wwuxl8rkBZ73wBoe+dn9rZEuJSETUY16RKcTyJmWF6I3abDu/Ih
alDkwQ+HNAVvATNoSADWgf/rM7L6/oOUaPT2TBcHrDCC8oRQ0v0MVAhsGFvECCqtORfBV6XsWu99
W3yvuNvAIistBIjxQ8ENoDjDTIWYSNV2DW269t1AcW/DP1AU/0rDg2qr8d0OrlqG+hNQp7PIZooN
nx1y4CVju01fMv0yQKj8wwNUwbnukgpEr83tFmnfYC0ZW/ROsLd3MIS7viV/v9Gev8T4nUYmfxI+
q3VVarwNtbbvJoIk7lJToCkqIdNn6hIcLsXv1CSvptHxIk0aeUqF9Bc9UaNT3Gh45zC3hM3d+4l0
In6ogkG4nJnXoxjKXkCYzmBTkNt/P6lJ82wPaYmhpvvThQN9eQVMC4pCQ3LkekCGyFklQK1ey1Xs
Uk7bPx+Vq1MYohLCI/r4dvVPMY/TBFM9iJsxzRW1l296x+H7ZqS5SKo6HGyAGK+n0pw8Ct0v1NE7
HFNyiRlT2xcfitFqvsiTZA2VcQJF+2ZYCrxnWQtlMtyJWYt+wwgGt/IFEYjGLgwzf8UuKWfyaB49
a830ry08LBCZf0lUzle7A1xU52e1mJF7iqfoQIzc7g49EYtu4SBxCr0XQGs+0d7rhh0egjUHTfGW
zxE1vKzi8WtfaHKUxSsJgg/ijk2mE5tWLtlq1pr7m4652NnkJu/E5z08Cy4X9NXf6ebPQfXy49z1
Qg5seqUFyW1EJaV5CL/hnb/v/Cqpsi6oVyp1uUzmsusbIR07SbQROKHN8Rw7p6atF7EnwnQGIKAa
WJ5VxPNwKO/4L4N8rsiZLWx0RczcPRdL8iPlcCaR7obhvBAPq/gi3Uu6Hd2EWldZtWv8YwBSX3Dr
sl29tn4QAD0E44rL8AsR7DOP6LsqcfAzYbAt0mHWEfCdwcUUtTxcm81NRfd89mRblYVw2XmZZUc6
mJYzsJ8gZRAJ+7Xa7LCDSW4APpQt8YszmvcJmsdyEeETLl3D9ghHsivfHmKFPMsZzFXlEA+rRO5E
aoJbeAvwGjbg3DwSxGyOeJg6tZVd8kBAJniDPWPAZkin3tpYuB2z+J0hysOeS3KhuOVKrBleCxgq
Ek/hswfSMQxElfySOupbEe/XQe+gN2prFgTVqBeEeiDEDnzG6UnkZfuMYkwb9QEwMQZMDm/zvX+U
4DfU70AyDN9FbIngPtzGXWHqzsM/xNlNVPF+tIfBhCIIr1gS5yBsdVlFqYPy9o0vH4O98TztPFE/
YzHRxtGNv6U8VgWeUa/1du0lsw0db0t4Gs59Pe1uP9wsfwLcoU6Jk3LfX41MG3GebY5dxoJ+YkkO
1IFdRt1S7aa5hHl4jMTQGNd8h5rZFL4GkaIiEUGKW2o5gU75JA0JXp97TFoDoESZ26cElP7sYy2H
PEvvx1QcFJEHCaUwSJdd3p3skzEgS9Jft7x9nqg7wmeUOMbdcp+JBvLefIsgzUypd9wIkFHPSi51
uiS6IQIy+Zn5cL6jFxvdGhkLONm+onJd3XfHfnoAvqye1kXFWwjJjmbdoxKmHzaIrvtII3zRbIlN
HHhhImbo3+KxCiV/sCR9kN2cqRkZArAn8A5xgVuk2sEFgkOdmV5tanbZIMY19ZirYy63RSoM4kvy
dIgN6+rIu4yDeosu9roMftw87R8vcIhsFQo4K4YlqWEqzRWhlq1owdX1C0hgfEsOv6yM6YRw5fTi
tW+eJ4bqma8TH65hj7OhK4qc4y2AjGsZ37FzcpAWIYc7aZK6hfEyz8XMF7ZEUuMiOH/QdzY7yPrQ
Mcd6dWujXLxqluX78FHe88Po2p0d1V1vC81WV3T758/c51iOAJVkX7kS+32N6+kyc/ofzsgNaozj
1AwKZ3azmERtj87dAyq9D68kbtLmAc56cys4IRA8/ZlpS7i+/skXs44Npqf1bspLYWfjYNzcYzjt
C2TEefd6rfx698O7/bsAXi64xil+queOpwgJaiXNBBeYB74SYdvXlere5q5lkSQr0T5gcDNtOH1O
614aWhok7vW5Y0KTTteftu7EEowqQew0jBAN013+1WpRddFOBfpFJWqIN+HB7ykVDW99PTV9vapz
iS3VxXgLOnHxRipfYt2nLbA5/bsaCwGjG4iJG/qOX/ull0u1Bd3UrwEukBUXUw+Ist+6dMUEdyPi
qzR7bVpdeXxmTTn3DWfcEtWafYNkJoV9oNcnLxNEAcSmyYyqg9HC9WI1FdxITNIQc/dv7aiMgzrI
jaGZPJqL4ko6bMyIrkTMdy+9gmukgA4dqdWpCBhx+I74xmcP3cKiUEtG/HaRdR7GQuy+8d6GgLIQ
DdsZe0s0wOfhT0tBg1MxGfJPvktiQ9d76Ia290Z+1XVEBC1o3mJYucI7VcyK4mk486kBRn8j0eQb
nkdA7PZpTgtESDWcRcKVVvzh6Eoz/aIjGt/ZPJC/O1BiwZ39iBbAxGAvAwdbffczmmXoOmliLriH
PcD+MPKAVw368x5lRuqShULSTPOzZ2oXEp/ZxwCFsVOQ+AcpcCA2GIX9ZljFOmgwmsYZEFAgzpKa
EXJOaC/S3tDDO2aFyux9XyNE21tGostt6MiQN0vpr41gYK4lrdKO2G80WWse+q/joXri4c6d5xIT
K0qNXAOGUfPTtHF4OIeLrnw/9YPJW1zBTOL4sq4fNzv6SlHKeFIpT1k/ZuMuP95R02xp9DB2J0Qd
d55jYxmz+fcBX5JvY9puakkKaAfGCdwrYGCddVsfVAj0o9ZJRNBoob2+RFlmBP38ftkocXA7YXcu
BBWnvzSEq50Frmd7F6F8F11Qkjd1E2WPLFNzVmWK53s0zEJk61JaSCXr73PVco91g92BT7nLI+ps
FanJF3NhXuP/LyDC+1bmpzBy11XyFeutbSD2ZBM2tYV7SQgAjpLjpbUu7blIkJKyzzYB6CTbBwQu
HYTnGLXeE9k0/s8luk2OSjzgTIt/kiROaLh19B1Fq+t5z2uIw84G8GbL/0BTlq8MgdyJywnte8Dq
eFHOOkSLzLMtrfImM8Q5mEW+L4xU4uEorIVK/BlEbkGxCWSAo3FxKTWOLa9KW7gBeELdqK7sSlI8
inyetXkUGV51jaEa4yG+7hp0O9S4vwO+ffbKnGz2EaVTWbOD8lOhj50l/jhRyDACCt3kuvoz8a2w
z+A2mRvSJsySKhxNVsCn5FkyB7SPsXCNlHSJ4W9yZfIWN+1Rc8AkTt6WVcWj4N4kC8p3q4Q3geD2
c7FaVZ9djDe5Ilad2XSD0m20V/VvgnouQwiszFlDAO07nCuoRVIEO9w13WeLVApbMqbQvkxPIqL1
O7VdPnIyEuNEsDVgGCWqx3s47gZWXuq3in49TcZgv5ffKHOOF7yP1dtuSkYs4iZ96dS+Fuw0PbeO
ZXcN5BKCbzPzb+hrbr8cnv1Ojva1I6ocfymYAK/OM3wtZjX7HThYGkhFb1E13uW6/D2lKABWM1TF
b7MDN/YzbWKm6c1ReSX5Q1rFYdfNzV1k2dwNvqOO2aDbaemuW1G8aedSgKWAI3w41hUTKcvJDLqS
8KBBfSWpbICXqTCcLIpzyOWJPjfnqVMB0ywmWbre3y4Xafu8mnHlKsVrNND0Y8SsyVPotmQ4l9/P
CT1OSyC7vPc/hJm/P9QupJyyVsoYR9mb9AmtX8b+4+BnJbK4lyyQbUJ1SrJuqBZwZ4pV5mFNlZt1
UueCoqGYw9D67AYRmDnnrParTt0kiqws8BSdsyekAcfoqNBAvKMe7KE9v6jawwY/QroU5Y3oycFk
VPWywnxojPY/w3q25Cuhm6WKf7sg37OS57oVbcBwpcLl/WGW/oijbZ4tTyAx7xM6BSHtGNKcsYkz
vzQdWpyP0jcK32rMOXfk72LOZ0rIJkZtq7qdSY/A86hFesuG+9zOmA0MZk77NqrP5nh8+IDXyAzu
CR1RLbVDwRk6GClWuOO3btwW5d3zBisdGKcYrMHhnzX8RIWaFOoJRApGhTz/wWWuukVAzJEl9umH
qm6k8712yhfsYyRQkRJJ9xoGHdesYoy++1X+guMi8JrG++mvz9O54fHQH9eZXVC83gO+eENEg4/y
S18UMZfhn9Iuh/uxIuI3xFagUF3VZe2w0jyS2SDFa1axyiFyDS5pn9IGlHlSD1HCLJB9JftTcxJD
IpUktMfbHrMAFXro15WtjjpgZAwoV95WtoAM4zDI1cv5guH0LyVtj93qpVEgXYRf0eztkMFpo2Hb
jb7X0mxx7eYrButSH5GIJu4J977IT43QBuZY97plHZBloIOasheIafRrrHVBhSYqGYGTwLT12buo
LIT9JYxASVBCoWtdMwM5xbNy1EktvQvPQfrOD7PluIRWoVUMyZZAHSc6uQNlVE15RNXDPrQZVFoN
ttahg77LCDrFvcUto1c2oTx2QrH8qbRw2rhi4v0xo2rwzwAvZXLKb5GCYtEmhV+itJCgrPOJ1kC+
BvYJXMLqXcvHc1hrq8ElS4C7nvl2GKoqoa4XVKJtDO5CDY+MWqLuEzYeOEC/TzRUat+givBJ8Rpy
K+vXk59alW/m+W/+zWP7fpOAfaNaDg7Y2EMahDe6Bs326+WW7dtDfdjAASB66aoFhUMf8lJA60t4
dhcCzZ3J1zpttVMYDY23StLV3AMfDKMoLb3SfHwinQgaco2ad/UFJW+o3GCX2wMdWCR0Ta4jXuSX
MFkHIel7JeP+XJxMZq+JuNU1pKQeRWA4OzRurHKN27Ma3U/R0XuxAXOj6vcKaEtv/7z63K5/W6jC
ZsSS9z6dZ74RFeZoyCzCsO3BKuBI+oTgjuoHMOSFvi+wlm/AxcM41rXFclYc0/Zzx/HP3ghdojcx
fVV5Lr2rQZ5KnIuFCrcZs4exd0Uyr6WkOLNPQrM/Shc7C6k1ZKTEQ0SnYWsYl4/4jMbFmd4zTT2R
NNXCnI7VcNemE8jAOLlR1w44Tuv7YwASj6tmpvbIhPZ+KPZ2xT41IuEhuFk+CSIzffDp4upcYRTJ
RzQgcIdCtUeo1RSLDuyO+BbCKZxmeqgMTFi1ILB82uz6KeAkn/ivtWxEIcXoUs1sP9UB8j5z324w
LhYPQQTIqFYi0EGfkB3MWzyCYZ9w1TIblaCw6qJ9w6/11aU7qzagpTuUQvOqe+nJqZ/UVs47jX68
Vz91cu4apJTp+r2mH3K/B2n0pJvrEAClspinK7vKvsOYr/twubiKfKdkPIVurd22gEywTv7r+tmq
EhZyobhCPsKiQU7M0sd5YKNr/ZlGfklbQS6KyBxgOwKHNYqiFfwsWmpWrhENcQXCX6NkPdERi9ZI
6hIHdw0ju1p22vDkdWHhdMJM8Gixkii6Gh5s2ysvivwImwSJumY8DDcycu+tk4y5r/med8RKTG3m
UOONzbcifnvul+2UyGTP0KHeoVq0Ltfh+8T6CDXEOE8b+45KYr30MBGKor8sNr8JWruu2QUK01Yz
vICLhaMlyeTBKAiiKDIdLumMF/JwMHPcjHQieZ7LaeAu1RQtJTVAEpNAONb839O2X/TxzYrWNG6K
8u1u1hkuLHYyQ0pahBcU1vGP/M5EPgQURE/lzPPEgz8VwiXtWmzNs7HdgNxIqWks/Mp80CgA89Ty
ZZEyHidO+6mxshGss45Wvzf/Lo131qIclAQDdwVu++6m4r8DIFrnf1mcuO/VgaNaX8DAkXmD1PLR
p2V6PxLmO4EqObo4H/o6TG7PfO8evEmpavIcHxHB7Gu3+CFMiZwgVlL+HuyvnySRqTGPpBiyzuAy
z15W+fLAWWfHnhzH+oVcKGwv2GCjew6+Jhf98AbBGzWpNbmRaXgbavQIVSmAjwa7e6MeiU5OCllh
Zbj5C067azrW5GOJYBBgXZb7XG7U2WF543ve3m6udAZ3TJ2NoaP2k25KFc3/IiZmukjNZPGBZoe6
TvbCSFI7GXOouI3kpAvNPfLGn5sX0EEgNNNHVlXdbvPg0IB9yiQwkk9art1CO6wbJkx4v3q/RqLu
cWrncbSCJE49a/fo3vZAj4pYSe++cnUKQRLVAOXdgzWV6QFdIsRsfNQpMuQn09q3zqPJvw72T79Z
zmfNT6NwZoBPQGVPxWLcW/q+1Fnj6JMDWaHhjymre96ZPDVb8PF4rcdta2b/rWtwo20sx+GfdZuE
+eNIhzsZ05dT0bbIqdZfcyoKdh8O+IPCofoLjtQSiy0R3nPbREpW0cIuwRGL+1TyrybsKSN3M6TW
u8/PAtnNtGRxqlh0VYUCGbvy0yJ/NZ2EWr1+PdF0mq+Pm0+TBOOsyfNueBqeJCb2kARio8pO4NX+
JabJP2Ts78H924jU9ANKWtaQh81I+4e9n+fi27L441Ygdkz84YcNRm/efoEpOZ2fw2YpEWxSPxQ9
rXqqkDsU/2c4vp/oo5kL1dXeSJQ8SRr+R9ic28Wf1gS0nsFNKOlpM8+P04NsD2ehbHVdjTM41KKC
THa3ezxZrIQRjAhUjekjuUXGQEqp+PHzC6iL/FK54kR28RV11FI8hmtaNtbR54aiCZCp6Y0k9zbU
DdmM0JxSBJu1vlZgC7w48t/BFQJzrDSd+u5APKQuruwVIE3euIgKM/9RVQt6BTntYZSex5ADwxWP
v39cr+1xjj7tXMKm5XKLOPwMx5JKMI4tS7L2anyK8ZCKNNd0ElLpLEfBG4JJGlBNqw0tJzLipEYh
bFZmsZMFQIG4v/pjJq+68JdECJpAsUF03t3agMambGkhmI109Uq/ZexeXHP2JOlGa7iJ+5cF/Fy9
etCUsx3z0X5GtslLNtsMKt1VJWGfbzgiEVRIxWOiLanVXv2khaCRHvyQzKn8vkDenLvd76m7TiIr
tIwrcF8vx47bZS6kxBmmEecfQdRhYpX8Zn7Z6fP3xJj77new0D2Lq/y0kmsTjLeMYb+gLk5bS8wd
BAgMvhyzkTwgxg2jFfXnds7vwDg/MTIYp6dplL3m8D4Q6S/11A7/0IZAdDTNeExU83+oDqrwCOaO
vSATa8vK2V7aQ67Qtk3AAfBPEwj87fGHwd24OxOXzvczkFuG7vehSfuaWBYZ7Az80u6H1XHEdKd3
Rmmnk6gqeg5EE6iQWJv8EOzDqNZT1GWHYORa4VLBR0/6HhtdI4paqthtRB8p24LdgytSyJStZjSz
+F+5crb9hEVcUskbxGoyi6nWlbwS+e6oyHMCGXbzxDZfbOg5GYoJtLltllP8zztuJUvIwAmfggX3
TwzKpk5v4o7PZQmi+lfMD6MIQR434UKRiPBNfmMJiob5mLBa/tHwqzmCs+EXQwtj+zbMSA/if7qL
6XQ5jbnKQIBfvWX9gYeRddmYUsq60UXFaw1MdW6w8GaqvPFO+3HTUWU+HtNgo3lwfSm28RNReAGi
Yeu99qpnlBXoDKbQpwY42yiZ7zRSDRYbKVi3bLsaK5hpNP3Q/y5koi6KvbKjqMkSh5aAdUzBQrBl
nrIOdq4lk8Wo38rpDRzvqkwGP/NqXp4ptlXa5TTJpH6lE3kHWEWxW6t6U4no+iPzYr6dm/kfmu/1
Itah6y7tIlM8eyiM4liINCE668amrY7NLnC/fE0nuZFYcU6ByBL+stTTPVnUwwHvCANc6beWyUnD
i+cZ0DqKiI1WPZVb2cNhAAK68qCPiWayVITpVTQhsyqWD2c4IdpZaxbNqoGYMT3kZa530DuHHW2a
wqnZTTD0MZTBMXjGcpby/riMmAOAkJNZX8YA74I/UKCWnjm5v0A3rRVSlBaQKqwrJwnuVueIivmy
tNhoWneYVUDw0ac5nkqPjUo0WsRDmPr98Au60v6xo/aTSrJJ+9Y2RMTa/jZWOzotCwK3/+LYcj9m
R93BYkQhc0fGLrNlm4JB2hVWH1HnHzji/UIUYhxDXlEZFRsGLbgGZXuwyPkT0x7aKbxaTFaiNoxH
5SC1fyxmw9UzuzUbcyofKbRFxg9baog9kvG1SW5TP2xcw9GdHYI6pQ2HUTpmN2RJv/UMInF9d15g
wsN1Aa0dmTWfzN4WWGjbgd6MHX/kXVjuhhiXjpK+Cno/KVu4dHLP71evLo68beEoI0sLro70DT0m
vjiq5972onToMZXvAaGBwxQN8x6llyNdKjliPv/3VhsA3QOxCKAecgxyDmsSlo8hIn9vT+nWFUAW
+f4QWfZ1LZ4e6OJIJXzowHrdIb05HmgaOsAJ7QojjVjDLkHdo938wZdYvsBhZ0+mExj0/QyBiALK
6Cn9HDBPlFfL4/WdFz+apgT6mCHUIKBqoviCDvHHzUb0SqrW3RK5EMNNvz6LlFtPnwvWhkajuCTb
w4UPYGYtvgWQyLALwwCYPk182VYMKv7vZ2YAm9hQhTzZcVqC5KkJ4JMxPw5tO8RoOKyxkIA4WCLQ
yH3L2jlcxj2ExGmbi311OrbylPs/if/6xl2+hoPu2xxTNtW98M3eR3US5gVAgxfX5/zLw134PsJq
SYCDhyPkAvjsVd/n70nXteuAdVS86SHuGfgyDkC99fhvX0eEtVN1ejk/f2pxDhfYL5u11CJaIFlS
52FonZzbt5PdyKgkFVomu3a9kRHgvJLUhGSAWexFHgN5C7REmDgaU9NrknzYN9gX2b6xkL5xZHfC
5oXWwdGYzrL0g022G0lsT5y87VwGy5cTH7PMRruniJdQWfxbur4oKg/BYD0Swq7Isih4RMCKh2wC
qdanrPKKxuGbg5z6I6FCW6a5J1obQosli5UEx1LJYuLhg97NkW9sza+Ve1wE4GdPDnUxp1x5iRjE
aSMD40PI2IWhWQjxQDlvBZ6hPHwinsTeO+9QxJOBTjV3OAkahDHnBmYxH9AVu4iYyRaan7UHhwiq
eA9Juz9RCTUoahA7foZLAkin/o9LlvovwsmJVjE1YxjmNYEiF0Y2so+MA1Eb1wvtWuaZcaRIa0/S
lBRbMEtk6G1MiwEb1IqDn8zZvvzr9LA8ar6JxY7cOb5eeyOzlXgh3D5WzyRyqPC6Kdm+35Czy1D5
sRl9b24LDIzgsouHs76VznypEqmv7b3sOgFOzAd8EcpqK9MzNeJXlwjcR0OwVTaQCm+MrQV2ycBY
FoJU1UvLYN4Z4ZdJEQvEsxfz0pa4yOQ9k8GjJgpVwNvuwWaVstHMzpGIEzpxO+f7tqsQHjRgE+Fp
g8gbrtvIRPMQCgoMUBnUzBzasxxon+jKgC6SRosCDUdFfbokVuy+9Nq/fzZbr5RyCtgcWCR4ynD3
jXUhEg1xstFgH6/5i3UilkLJmNM+DqXVPpJ2mRwrjvhT5ZveheuJLe7ROvhz2N9Ji9NIO+Eobi/m
3bDZ1SAlUvkO/G2551ctV7VfecgnNkoeSxEeXOZbN9sk7QyQusazT9IeHeMu80Pjten4meaZgKbq
d5/6jcrw0sRsJLn1l8/aFkDVUQ4h/E8wYsgeCRKsMYTCQyqYfjfvBOBPYL9UbXip91VOrHkiK9WZ
5hRVAoeu7C+3TmtxDzuYPWB3L2SED4Tq7Jjj09VQJcvSDoKwQ5o/APHceMw6vwJMU8pDbGva0wNm
CbsDBbr8CAxZfUZzlPbQDD7Uz/DBAmmVZDdT65MmWuMnOCyGbFKxJ3qCOKV4beVZfkgr7fqn60Hr
xekVBSN2hWMHoFuWIUHpnwBWlLYNE3djyLI8zXsy1Ur4kZzeg4tQYQFa7TFD4wnj1hzRgTg+TxEC
lOfr+bRFi4PndA379wTPOjcl30CHCOWfzlnftM5hJQ6pGN9YDRgq0ZjvAaD3QG+OsfXVd+lIUB5D
KkvlFe5xxQQ9rvFEFYcDLiE9DaslpsSvz303GQvdisHGuLm+FAZoUHqBDpebY5Ff27hRdZVGaYp3
dEhK/6NpkT6SNStzNr626FdLLhJeFFTrlD9cv+zfdf91NhEAxYg2EvNvxAX1gY4Y0AKQQyaCOAw4
f5m8Af1BsaheeI/7najs3fFYiyZiTgbgc0PLy3C75aZzPjbGeu4dqS3BLmKPXpnWgsIV9PWN15Oq
j8j/2pzwC508twj/X+dO9yT2UMhfEwuOMNTlEprC5J5SDI8gMtSfzkNK9njlyXp8M8oI/Xz0WA+s
3tsxP0Fw5/CjnVyL2cfpZN6J0A+p2RTtW8dT0feINxzi0u4N76BxHH6xl7QCPhDyEakorIZXDSKS
dhItRtrWzo55CtPlXAQ8bfluPgf00qhMf/N0Fe7xUg2shOAZDt0mAt/nUYK/qBYegqqFWQhLwrc0
fpnccF+M7R9mb0Ny8W1loA2brT3WBBsbrwPCYkgEWly2CkVHly8VMQWLDjm1cvG3e53Wtc2KwSUU
pDFd7ZAOgy5XMhNz4HapUO+FgNEW8NK58dOw/ElM/l5CNC08+pU/IjcyMDBRQsNzZ+UEIvh/rMxf
TYKb+Rupj9IQie7L862JhCRpOhDe8tedIeFybGORdAwig3as4jOE6ajDf+ISYmhjVxLyXzJc7Xzy
ceXBmh/xoYHVkgXJbllTz6UhXjFZ0PkhelGJKt/hHGm7qCiQLYfPjViDyMilEji//S0vpE53xxLW
1g62XnE93LSiY9PGedsbLoQYUxR7ZuBxA76FiAbfLoFJU+AD03x9/BwWrjst+DjSmhfSVi8244Qh
DusOPHVzDtBcpLO8ZSpN+b9LfNqr+yPmU1kQYBaR+l7Zt+3Zu3smF4JppRRzTv5ufFXJg3ktbWJ+
eB9rqYvqWU4w45TKzUdmLRXvAbEZDlGmWIB0B/mDNAYDKtWRyFzv2Mq000LithFY1XHIOnnkPkic
0fSFlGsA51zL7uBYS+Vu8W0WDysDA5K+68Hg/Ox/v5ggLQoOi/kNQRz1sfMaIP+F7uei9tQR3yRw
2alIE5YUKGU1Dhz6RC8cL6vna118jDhOTHNu9ch4Ao2JGZeR+0MRcX9GRP00GNhu0mVEgjoXyYbd
/uTGtbXbZ2f3r9TJ6ppqBncInnRDHu5/+bHxNHb8Bfs6AGAHih5rXObSDUHx3yWkesQCEM6sa216
Do29lYPtiuxHpT5hTGJbwZq0kBPtKWF3a5JSGTCf+98XkKQE+53YuuFZ0nz4I2USaC8TQlvesSu/
2bthOaIaD6xgQisg2+EJdUyefCbgJQbLiLMQG5FJYm+u6DIgX4xeMNGMuyy275P4jhDvzgrwpQW1
x+CanTLKyJlWYJcDlu9wEsKkXJq0uGrO1WlK03B0N1vP/P1ypp9JaZYK9qiSu+JDrd0hucYnWBOC
LztJooYsxFOyw6UQrhn3XcL5Xc/SkrJEAyO7IaNdm1ZNOET71wShvIwlDr15AGPjvLONCASkGKax
H+9FBabXVyG8tOawGjuR5D4evR8SXfc9hOS38i+l/luS5r1KPm49wRTJXd81uX/JZ6CAfZX7uvyD
leCK7C6bSXU3Rso4dqhtKy7QlQA1HoM/HgZ+g463mavlWf4EaThCQsqba9DtM+9UHBJ4u2J4iRcv
Mzrvul8aSJyC9tb5Y8LkMir9fEqZRxt7yfEqWIsrW5NWB2S7UAScuLrBB/G+QHwtSJGUdNpuedrQ
786bXTzoMUB4o02W2CdFwEbD3szxiabx8QxBlWk7YIZRlaqbrEulqGvwbQQ4+wmUFwnGmwPxhW2n
tk9vR8OoGjJoM/gSeIKlHrnI2WzJmp84o1hoJh705/YWOxaF8VD6x1Fo7nHW1VpqD6+TPsOhf7FH
V6h1eml2o5uXZNZZfmNFoSRm91f8kp1yKYMR8Y0O9NNekgQUhyDdc1H5G3VxIIzj9RKIjgyLXym+
nKgdAWfoNMX+IQuxVO3OUeihtSeST5sqVu1CAzJkeq6W1TMPwQemz1qVHfPJ7hO3I+G/uMAh4vq8
lDIqW9hdPyKXxu5u5Z9dHN+zNvKkOy3V8o/QEbj855kJi+AApuiuY4uiLQCWPQQprEpxca1+do/h
A+S07wlfP0rkCdfcoSbTi6cQOpKQ34s9Wl9q9GKRvSImOMT9Vf6vJgdTeJ4DRLoIFYULslAy9tUs
cUylr2iFii3mqAruYC7i1eDWfKJpV7Ufcawb8VwovGy76qBF/qHLBJGajtHNCPjcgOYG/gDrlSLZ
9AlHROXdI0kbVB5+xYQHL6Wmtv6j/JcA5goL7IyjrL2lhH87DuEvkWFj9nktH9qtbG1TExsmLJYo
YJyHIJPgQdmiBbbLIVFpa0QzpV3atHCaVytEXYAsZo+UOVgM6bzlW2eAagj/OT5+dtZke+yHyKK4
rxsZ92Y3WIi8AqsmZb98rLnOjiuee0YCRBzEvaH72VOcE6AtGJ2GC/bs5cVQqThNN95NAonld6FX
/kwcYBrlxcanRef2jBRecLxjs9C+6kL6IHv1IgzV+vKkp/4sleiiJQ9FkrVNLHOfC24qAtAXVAKP
jiQn9TZyCjE85XtmS/R6mrbzeMBJFVDR9iQ9SvugnCdcjcnwlWfsWn2T22B81FHAFlkT2jVt9rm4
Auu4qfX+LEWWyGDRDwXzo572W/3ooHO48cSu/Hz0KJlNVQdiQOkeUvXJT2FXjrh/53nOntup5V2G
pxQLboImWj4lvlQO65zwt3kLA8y/22S0IyiYVpbEWqrFhV0h3EkwvxCjlIajgubWE21gxj7eVnlv
4pGY8Y+a2imHFU0JEfl3XRUlm36bMO6ElW/9igotMJCIQCnss0DEEJRk1IrogFsbx7YenWzKAGLJ
7e+bp4KQyoJwJRkVr+TSY4udYAWu6fDhkDe5G1kq1bTlk0rlCpEuXNOKM1ndpMRokzSUVk7UYWQ2
dtZhJaFhRJv9EbSQO1JRLK+CBcJUXxsFR4BIT+KGIJbcQeZrR5em/nWXw/9t1Sium5eXruqZHE6u
1ZumpC10ufKeR7AFLFbTeiL4nEhnesMWmQ2WbTrl8iUL0c3vee7SVIuyNPjno6HuAeAd8WkVHObg
rwl0tk2m7w1oXriB/kotfQEk1jintlmoT9t2gUAv+s2LBF9R/NhDUTiCTDu7zM6LNGbZtyzucBA0
VIJfugDFiU7T1b/BlvW0nP6+Cl1EmsVoBwdidrSGIWvd1lxzETt47kks2L2p7av9jigfTxMq3MIe
wZLY4cQc42w15fnKxLK8Zsqx6TIa3GeR2NHKm27LN4lz/jxuuKDafPqekL2b07UxOh8TxqVqfKHb
Y3kksre67EDODe7TSwi3FHBur9UP2LpgiT/cri+OLa0+bsNiH4lYYy6jcdi7oViumitJ+2TM9dBy
6JIpVCjyn1yIP3MjykX6SnRYIT7gY4HzfiM904ZjvjN3yfaO7jSap/krB6xZt/6pj7Pn5/UzD863
nZ7IrINs9DHs+fD5kS3SmM7agbfG6XlVZzdE8lRcib+Z69/e31amS6DvAkjbV8GHYVaeFGHqR4fA
GAQB4URNEfr3IZKmsSESFnrKcMrUHQ8eBsfIrJa+zB3awInmYCiCDn7QM73oFn+BZd/owYYZ1cvE
DbmIJ7ENQTQ0yHoldW1g93hIwXT0/ex2tCifUVsAMln23ZrpEtUkfzCZpRTT1OrcSM97ku3gtWe2
0/M8gBDcAIpXO6RzARJcXrebWDa3An6Q5fYyC+isKbzFR/Z3c/Y8+xTpuqmngAJrI7Z+H7oNRvwJ
/VJrN+wisA247+yISl5WJxDHQ9jT3HLPvg1SQHX0qroeRYrbYkBPVDesi9Y3XThs3cZdZobsPB5i
NDzTrBecvm99Z9e/4xMsUNz+kxv4haMNWC0cCV8itFWpmMSsYPifr6wlX9LO9xw1b8VPKu9R5rk8
PEbw6+ejA7dQLvFKRi3xsDhti3kBYz8XdgeQC0mov95QzJuz/bq7MZ1C9z38UpDxeSC3ZE3PbUjQ
xqPGhM/77KbNFb1TBgQNcbehakRujgnv0j4giYMYUATycK07vfSMqssWllLyz4tAduahWZLXTPgj
186Yv7xd52VUxU8yZN2Kh8E5FTqmB+ch3fcnOxqMcbm7rx20VYF/B3vrnw5xkd5oGohGcn3Ix5MB
4h6IMs4GqFdhThQlMlOzy6ZMaBR9veGIsz6al/PHOnNPj2H6cyxeJ5wsRmtDP3sQOEiOBfOGHLMK
LGiFg3aKso7axETVhc1kuG/GfA4r8XTFsrwHJy6IUaFrY/nQzPAv6Itt5Sao6+I6t3aQQFcsGJDv
kXkyAo7LtmLZKEKoOJuUizxN+/vZKVl4ttvQkO/iN9MimVnXSfWEdgnprCPjhczZTNtZnBXOHxQq
m6HY2Msn46cm7RJMnAoM68u1QvhzPJlNGcPTQK8DMfGcXpP75i2RbhbXLqPe8/Q+MmNW8dA9JNlL
N0phDKwI/hD3x7r7nPtx5cyaoFsUhsJbmzHO8K0McUh1VNsqrbWztEziLf1vmCdQ/MzkF2omjhmt
HcPIm65Z6Up1GKNqEuD+2OPBpugVny/QaINWrS5Cp6OvkdNZ+D4iRrkcaVyojhp/lPUNTgUvsrMG
88Hj6WGqa6Y36OThrkfS+gFwVtXVBlMj9RMzn2J0xgxw9uSn+c63JxP4SWeHNgZnAG0b2ty29ZJy
y1tN73u3iOoo+blBN2I3eEQ63m8eu8uwj1TI10AkRrI0jgHkC3O41SlJdqSdXHM3Zdyg4DNXTQhU
cIYzg+3Q6LmJ3PMrp1+Mym/Izh3R7bdZPHsC1XALbWbO0sftz3V3e11Us8zP5tCRtBw3G19MvOmL
XgkiW0MSmh0tPr59kdGZeGizGMwo34HQGNXdhybnaJO7mac2Mi8dMn8yVQOGlsm72O/QR1rGlp7W
2R79sXN3gqyIhPQCPVnTr9c1RH/TzYuVpO86u4h2pRLlOK3NZvcRFmv0AcaNh2m2MSow6cfqFv53
MMCiKq4kq0NEPD4NgrgA/iyGbEOlbWfG3oYaFX83WmJwq2I9pGc+n/bQDoButH3UQfI+CGqbaTt2
/W3CJuLwvYOg8/x2QnfbMgtBEyLMHYP8EFIBzUK7eWWE1qhPtwtehGHNKjPhY+BmzwkQFni3bFgG
NxsAUJdEtFdebKML/e8sJpSNUKFz4mdsjrqo0ewU036iDCsKlbMU/vY1beZ3jjWB0tHGT37lGcIO
xfZfSwOkItYFzkedkAecZozYT94ZOXaroKr8bCjSu0TwW9P+//xlpZb7yyqxxRtJBiZgbXpcsz+b
fVSlsrhjhETDVl09EIFf8KeraWn7/18LRzljOqEOBQ5f8dDgxB0/rDswKcM1NLT4lWbAOAkg5RvD
A8OGzioiRH+K7F2Nui7DsLs+M3JMGxBitaypLtG34FHYUCO5PlItVHHW05AdyHtT9K3IBm+AIhwR
0+Y41KcwmC/Bgz4XiwIdMHAZ7AdeteyFjlDg/oOvzriCLkuZXtEexpF1MWIPqThfZ4fv4Xk7zhKR
+mkldpKKNbInxp1+XhkZ1K/pzqrthuiYvfHxtX8GFursxen6FbLfcBKwbY+AnMot9PxBTUR9wQ5h
UiiVBOpanukMJci52kE/3LKt7XGY0GJkzrmifzf8n6GMmsv9YjL/fxSNzgc0f51P6Z4Xt4cpUZid
/yTzScymvkNZuQhbJn38wxJt88QwoCLXgzyUhjGEfkgoazNbURDYljdHDCcAS+BYCrkaGZIPlgoG
8mmVV01otcvjmCu81N8Czdmrwr7zB9DF43XAOhld0JAAOkAbpWCPHdD30eEbg3SqWGIbNi9cTki5
q34T+rV7A94e4bOSuL/UbAELJefJT8aq6BD8tx23EDH/u2emX16WKhk8/VZyHcFV6R6zmi0s9HMw
bGUe0o+2PePPFsN/KtHdY6UwryS29r6+Ttz9GJVTmVSWkDgyyomFngdKOuwoKBuy7tTz32K7jmxR
09GRu4fiSWSxBvOdQJ8+2dloLvXBvymYvpvq6Jo1FqNNPhAdHAicha0W+soklznnAUx0j2XO0adT
HLF7yy8AwJaPd9vC67bofkJNN5wLmI/9BvxjbW15Sg+BzFHONfo0687IU/wT63M61tj/1EHJu+fg
hcAkbDMo2GUeVNioyxfqr5wPr9CHkm04toovTgq9LP1WOAQAEzXy+X8AlE23dbPH/NJbTKTFYDmL
Kc8b0TW+dzQciO9ntqAyhYMSnEs4BKtEf/PhfySb/IJNkRe3Nnza0DeN7jQKVq6l23Ml1tQlOaVJ
6SYEQkLq7RwjpJVbLV+iD3dMgU2ImQuhzuZgiCTv2qKM31B7FMQlvF2m4RYKE3qB7E2jeSzh44Bo
2sNDBc5BM9yEn2NgJriWL2FEVna0JiI9wUvHOquDHsmRtGMOOu6e/VCePh59q9oNRh0OlKqHoKmr
CGafA9DVF6Mm8+r/nMA9qwN/8TRW4kUUh0qHRN2IXJY3PFX/DE7Ja+wV53imr4BuWmFLmgB52frA
EltEd+FlU6xSsfZiDrN+hQN+gL6yQsJ6iJjqW/pHWtY4MVlhfArZH8UB6v1ouXjaRz7+rvNj/CjK
oRdmuCtWE4JSFORs64QIsR3Uspp7bNWkuvJZEuvsTFCq6N/WqeDhPS8TtnVCN/gEJIc/js/yre8u
r3B6NIL8VsCJbhpOI1XBFlvHuqL3KpGoCUXuxexVzcMCdJ1r7aAcNAS7v9BkzZrFbMyWI+IaMxUd
DjOO4It0UE0OFG6TKUBINh0di+QI0q6kB8NENMdh5PtUCAPfAmo1hSZHdFbpQht1IAMbpjfY1eSX
sYtUJoPc64Yjcctji0ZzT4yz85qXS8X3a58Za0bv/Oay0UV9UV/uaL42SX7vsa6DtBg8PBfoCsyE
tRw9/R0tGDaHoWwvj/JTpGYSLRSuet+MTAlpyPyAQgBHA/T8t/Di0K4/8gCo4CbQDkLfiXrMSiiM
xI7IuVvkvrD2CmjhsugpMyJRgJX1T17EOVoXMSgSc/IgC2ZCAfCO4jN5AJ8QKbmFjspPomU2UhVW
DxC8icDBOdxSSmYzeUIdIYnrCm09PqESUYoBbxKcqHb4d/BILqQAbB5fgsy6OABLe51ERx3MJ4wZ
iUwbQMpOtwENrtt5X7KyiRPO97ATPG0LwCqhZMMUL3knRClA3Y0qXvSvAwUFW0cJDHJsMcr1Hnat
6cn8P4rAGAbOP/VaZvnnrX7e5RXuB4HXanLWzMhr8cd1PMdm0+IDLBVIslENQu/YmU+u7oc+BLmP
fkcDep9vUz+9eavAVPCw/AiRRnKJxIQL5T4dYE661O7jluTxH62ArtvItWT8shDD0zKxJHSHPvPo
W4RI5NqO9M9rxP3AUkmEWmfbkDOLX1qie05zKVSwBQh+untB8ksOjaZqupPXihxZGt1qc6lYTnO3
nQzAAKLIUEZ1H4iLgAWd3yqj5DvCLLPKdHupQFZfgSQBoGe2nI3NV5Fup+Z4umlY69zWKC8M34Kz
uW9uONGSreNIKspd9OT9sc4LCnRMyIPN1Xj4xq0CMzyd90HwVG/Oq8ispTq7wpsEVTXsztWMemHI
pisH/GGNyfMAeyfkoLDFPQ6kIK1M+eDyf5tSjNEi0A+ws80+xb5RDc/01js3cQZPy4y7YoLI7AAY
XibvQhJabIm+KHHxM49dKP1j1ULyfDDLSDDwgYAaTxekxzzmLASwY5OFhRkf2wsrzGIlvrULQK6S
vWILNfsyWH1oKXjYCXwQWo/kgaYgZ4Rz7JJgRVn0NOsDegqhD0CnvPPSUJgOWZD/x7tAKmT56IH3
s8s0UivrgZHBGgS81YV24xqZ8zSzQ2Yf+T53mWcAnC/W3PKPg8Md4oTfktdTH6w36JhzfL+BR1BV
ADs4RnX9V4rlj7bbsZYZKvEp+mOm3RfXYj6VBQeD3Qabcka+dSuZ1kGMSEEAtxBvjjMBi01KGDUS
vMBNt0UgMFdCdYQdGsrd2lXg24F01VEsjO32F7eVynzsq/enhPE/NytdFb0BoyTFegGj/L461/zY
c+U8ZRQdFjL1+K/NP0rqZ9tBFYC74l6dbdJoK4lOIW5vDX7ZXpYt6qTuaxG3rXdZW/tZPBgmAvTk
syuUMkSXsD6isRJCNS/wvj4Ikn7YeOTy5ATtgz4Lpg5KAHScIyP43yWgJcNdiCXp9nmzk2mQBteS
vGmpd3LNFCihDBuhpwv5QG+nE9S4nTlwsHpO2+wbabfQt4gRnGGB3sYVs3fz/RRby5Se0COpmOrl
PhuNYliYyisyf+YWvfsObAH74DCOfV8AhHJktShqD32ToYZ61oSDDwwK/YBm/ldy/ZS6kj6SlTnL
yFKSHM+e4CJh5vGr5GdlRKbSSp8i1kkXSKB+WcriTi/UuhBU8yPY87e+k05qDTpqSTqSQ3JErLXX
SmpK75urM8VAVOdDxsFtQainDjuJKGJ5b1PDiGXS6KmpMvBwgzlRpvSh7IXQHbUkmHIW79v3banU
X+qgvR8zvIkyE9pua7AF9iUuHHcfsWQ3l3H7v7KPJwcIiebb6uHODoVj3HfdZBuCZ8FAMLu4e7bg
itVyNVKwIfVfFFfZ9GvbjSts0GgEdM0DBV6FcqvNCX9P0Cbzwm13e+om6MV2g3Yhx/VMOizNPRE0
RGJeeoTcRhUATcQxcjQ1sXEYcQDipSBMV3YW8/SxVdNkQQdlMS4NtLJtGCZtjb1kmwL+81dBXz3C
dNztq/Jvk/nW9F8wB4ZLyGrzwzZ5ugYdt9YSVF4G6r+qHRRFRhtSTgz9b/pZgufaPFOL4BARn8xT
w4tjjIB5wqY0o0GC4MXRDuLhiQ9sOtGx5ZNVAlrZFNUIWs1/Dv60de/sok75TtVy1+Pe3UKYEIi1
ccjvwjEr0IJQXBZiIOs1VBf6BZnE1+nq1riNWzWS1EQ7sql5S0ENYuyLoHiCDZIOkO3HRsPU+jKh
TDiEmQw9OUKmYgi9+JpIOlSocoS910+J6Fx8Xe7qxMOwSfLDyVx2hz3Vwul9Cj0zX27r/1WgQkG/
kwtnZJfcLVKFgZ9D0BnwT3QUEhEHFxgI92cAVnRwzJwfp565L/MdPYpMo5XZcYN+haFCOXFDxgTb
jh/61Yj9rh8WEDWVHMOY0ZiMQFqZzuFICyovylAZXVPpNOraKOBUZd641q2g/HqG3/KA79t4AH2r
h/oEG0BP9CQjzkZeH0vndvSt9WoO0taWfOeKeWaFfVTril/WsAafpsTt/gOgcOMrFrGqil/soodk
thur2pI00dswTyZqV8AO9J1Mbhr/+wP8L0y2TFsDeJLX0dS0+CYr7+nBUIe5AlOjtbWo0Je0U5Dt
4mZrKY0I0HOn2ayjOnH9jsW6vwX2nquFUUTpP3xLvjymbX/vvOiLtOpFN4dIQTkS0S729pCENKbx
vbbdT3j9wHJerov3YKjLZ/UA3G4/Jz382QFDu0ShKlOvi7hU8Ghx/1RgOyREW1xVD28yqddRuXDZ
2RIHHu5TrHkyDzfBUe12zjhSALRAw3uGFoMXcmttRmU5vlgch7ARp8b3DT8TF7dPT3IYD8MLtPNK
80xubcnmRFxnfM76C/SIi4bCQHrDiyjfivLVAJIVL9KeD/DolXIDI1A1X11XMFRcUsQKkRJa8de4
Zj9NcJZW4Az4GApHK+X19kLlmasLQCzoPE3Yvao4EcALgTy8ZHmVn310EiLpFXvZKgbPeBZW6BHw
Gfgd1tdFihIuhO+/HV6/n+TTNk7BtV/RIuAB6PFB6YIDC+usDhkmTKyarggr33Y1bT2uOimlTvd/
N/E/Mn1zRJs+Dc7WQR0u0drx7NPVj8U1d+whOw1SGMMz7gO67WljCrBrO4Oa76dOybRv9rJjzRBO
nOqmk4qL5IKQQEj26/jjkstvqyfKh/Ja95cNEtLrLJZLNwMN0uGFGRq188CLlRGB1tUThWqWi8O3
BPQNmcu5U5DioeriRWb4tIH4E4f4H3lpS7N4/3r0CEaayvXlbqaU6ccEQplMrXpDowiX30K4YKbB
l+KqnW/EuVxU4Ab+hGOJNKQItjECoZaLYCMfbCmtOxYCWfbmy7A7yo9ov0Z5ySBZX68PA9OaqWbm
6VHzEv/7go4XiqjiOV5LvZF8KsjdkrZF0+INjO/xwmtLsJdid9ZEcsG6NbkARqVVoudIxY0Jg500
c9U+LNRNU118mQRgV+ELhHMCxhDEzzemnhDyQXPFmWcDj+STjljUnDBFVCC8scd/h3b06vuwOd5B
+qOr20xSBW3vqGFwMIMpr0NqSyL4KTLYJQtgvfFnBB1eYAa6EEzNR+PGiYvaCh5Ed+vh7/39TquU
VATaT6B4spNZTypeomwFa+CrW6OIKdtWRiAL+P6fhpT43EHIpajO3kaYArbVZfwU2Uhi8X3kopCu
IbL1G9L+J/nnRkC586tYzS3oXTxpFRo86AoyH/ate3mPrz8eLeDx6APfH7yer5D4VT4YLg3ataTY
l/75Ny/hDTGq6GmYVAbC5iSCTzXXirqEuHu0nGZfKtopNC7BuNxx8jdzXMfZsllunjqDt4/kOozz
5UaQb6CHtvLdYyvERagbegescwwbHGMfIemhmTO7jsg66ASmyXWnNcdO3WgepqT7S06sIbTPF1n3
VQ+Lnt6Lzl38zp+7se5oZ6GdfrXweMwUgyQertMjj3yNlSdkk4L6tt5hBs0MsLeyfzoHQE92JgiV
zax6GjoKhN2V3lCxeELoO08hndHLUtGCKGvGt1XK2w7/If0iJco1mLt1FCzlt9KluLJGzWo8q+DB
2x8yW8ggogh3ct1yF5z55keWclg6zrH6TIrj9BTO3Hw1CFfKUme8DhLwEmEoDKkD6fHK44WU7Bur
ehSIokROAJ2fD2kQD5e74lddNRc+ytXagsN0jEWtd3QY4BrUhvQGs6f2gyRWaCYkg26Nx3t9QGKU
PZnz+uX+1mur7nzhB00uYrbUBF1A0pN0Jayu/pSQItCyFeKvFc7tRt2xAAInc/eaH7M1it3OrO6z
0NjPZll6ItxiyqRyx+HzsUCaZZQASLRyEusBlJm7uesZlgDAn6RV5rlB5VoBLo/AiU5JwwQ5oFPt
qTjctRqMzttdcOxlK28iAOfexxo8+V6r1ncsLiNXQWndfv267NoOp1Wfb3jnLzglirkEQTacwMyR
1TZDE68tkjhta6CPXn8LHM9TVXUJkPtVe1T7IuXe5c1LxdihMUgdJrkaX1//6th9E7/l10JwU3qA
Yv4m/agblvH/9ehNxCbio7YMOBKGYwLjq/emZMrJRQEHP6eZ/GmyiuZPo8JG6Y+MoQT2x0DZKXAs
e2lvdpq3hNMft0ODetFXJTpABoHQ74I0LoCbW2v/1JBdkHJNh7et0C/V+zvV88/5E7C9CZ0ThJ42
bS8+CyoH6HuuG6FCOu0CwCEpUy7oA1eE2Kg4K0lgYnjMRRu0JGL5IENU2I5rxRexPgP3AzMs3lT3
ts1MOw1GwVghyMrGu/8HwbPcQz+zgIXXjPCB78tNm3T5Yzo9kR6g9YSVo+RcuNZrM24EqzapTJEh
ZNNnMH86sIcjs//txZ5S8gUNLaVqSJOpIwW5qRrx4cmk7ORrjdN54mtND3Gx4b9zn5qCjpfQvXVv
EhRHi86GB2q0y4h2zDHFZ0NQFw3EwQ/IDV5DPpSDegVbIJaHnuqJgifNXchJ/VwAQuIuVyPt0rrh
5RD7BQ2YDMT6NOtDuV5RLQltaXIH4ccFtvXmZH/sHQwpsPkcXT+EmL2FTSahXC+Ly2oplcwSRaOV
uAhAMXW54R4zGx8/vzCCCcz28/tlUcwukdX0x0NY9oy6kvGVyP/qIh6caair1TkgRJui2B1xKPA6
GZ+SUlN+0BGt7khwWrRwfomKAT+1L2wioh0ly1o11wnc5k9GyE3Lg7ha6hBe/vPhO0/xt4+KPv6i
sWlTCkDbbxERrfJPwbt8kErLjETjWuSo4JhZG6jYNHYHwggeaxyoJKd4warbx2kD05IpBNgQdGIM
JsaXX5hZ5ez+94bGUJpBGPYxcPYDqGqlIOJT65whj/dytCuABk9JQAvWSbxdg5nE2pvwn2AZ0UO8
sxqTvr5X1wt1jz7R56JSIDDSFOrjlu6Lhhs5FlL5ePqsFDQ348lw4k7tQ1crPDWxoxl5dVD1CZzW
VdTWo9GflJ3fHGv99z21l+W9ZkUup6cdgqNidWSxg7X97hK4KH4YeZsPlRjI0AHK4gbY5/lcz+ZO
nIhcq4k2Fx/c6szKflYF5lqBiYTW/vEOItHQe4fDwGElGSdginvsBBY7LqkBSJndNNpQwAF+/YD7
xN5kEZ5Pfgq10iQwV0/A3B9M8sXcNDHfmfzR54BBjLKu/34bRwChNlh/To57cZc75qkAp4ikse/N
JqEl53tvG7p7v9XIpkAfre2CagWSWGFJU7GENUkFGLpRjMDsHNwv+lCNaA8DG/SYGVZ+Dw0RuND5
qmFDlhHTWGTy32AZeQTP7UC1jV9B9SPa7Fwhdd2wxVTK/JBmEDoN6S2FbbpEra9Il/GAB5gHWjaF
tGDBHqIcA6O1xPTWGM8FVpaRnzuNczVQy4U0MIgM9H4RJv5P6lU3HNaPm6K6HaFeYd00gyoxEUib
XGU25ZFO+QcHviFEWOtwVkcoLxk+rdu+KCh5B+B2wme+hfQC2mlf6S1h2picOokavvhnmESBjHib
y6gyd1xJnYXvTVQCuTZ7paN0xDEwuSsivseehN55YZUD3Lmg51w4MSWolIjD+TKtDBfNeL7TqbfE
aMf9kGhNyQkq/5Woougpd+A/DgQSMtcfMyn2pDHNQ4TRR6B6DUDa/YSx6WmomBlK1SyohioCoZU2
FTwsQH/Lo6SB02vMBrS49Wpa+Uwx4/GtvGEmal7WSWUSUsu29grkCwpC+audmK9f8ke9j5b8ftoH
zgxqyxpuP5MWu9RNL8CgSYnLSn+Fjq1HZLYe5sn2wrW5Iku5drE6I9etRRHthNT/+q7f+gqyW/T4
3Pq2ZxhRkOvyx3+PpYct4y6DUJv2XmaS4jPvpbaFYslWMb4MF1tmNb9GBKvC1n1QW8+rVUDptZwN
lMKaVX4FwHu9+zgopsJOg68hoJ4L42CoJBJpSWhe52HAa7iaPTK4vbLHqQMPuS7nrV2fW0piNUNJ
+LUIQChjGgrTQevhAw5vBM+WEUJNebHuGDNSisRHa8tNSdjBDNEoFXCXfYEqhrwTvXyQ2PnUpKI3
b354EMs1rT97kdlxzfPsZj5JU+GtsagsUIv7kBTC3c0lhae5NdnfIPm4a36qhofbIA2je6GRV9P+
UNOO/wNzp7/R/V55v2qXcRxKcdJdi+Pi8UfvF6h0oEmp6lITVoP+oFbSBu14AbhPD0TZMFLZsQKH
eA/2AhqWogV6IrB8gWgOw4SVH0VTmNZ4FBI9if4B/tYIXaOSDWyq6W6HdMknNxnFWVXUT8EdNFcn
zqOYp17lNCAFN3xKzozyOHeVlkQqmH7h+ITwZAtq/acCFeaMcOHjBzaQ3YzRwlAqrBYouBcKwzo7
whcPNvmhMFQHLpNvSaGVjFwATsxSxkX/9rxLwLkLqmvhd+SO8CjLfXf46YtBVvu3N7s03KTWpz+8
wHmgF/TqQnh/NKcvHoMThc5wD2L5s+qBrkDaveeJ2T5BR1MtG4geAmydmc8gEfUvgT91Z5viLrUV
7Ouuv7A96g1r+0O72nTuE636ciqiUez9gcQQuaSpbHvRevFxmtuGuL3xCBBfYaartkTX2wq83W72
uPlCpg46vjf1dTczAf9Xdh9kyPFuZUaKPWOh19aP2v7gVUKgYBIfPyFkRopAcEpHTA9ihdnpnyDg
Z0/7S8JvsRaBpQwEfWp3EdFFA7wstxhpQ2QwY7FyXAFmtVwxdN7g9e4YqBvowh3nMY/Yhk1jCuNs
uHHxFEycASS2b2pTEXsyR7TjLy0TjYdZeou1ifIhP23r27KtCS+JQfmsRB3TxCemkHIX94tyPz28
aZ9n+8BD4JO6re5CdJALNKxzdl10qL7fo+FscLdgzTIUnExp02w//YZg/fDK1sf94aeDL8xNIc6D
It0tWF0V0PIxfJWAmlhdJN7kNQHBiEbPFDB0veEKV7kheUIgF6cnmgqKzQpybtNwGQIRjRUvks2Q
u9wfaF2OcE0MJ6OrLCPR65Pw5odzfCArwj+SlXw2y1ElaNKpV/+5wZ/ls5ILs8m+wnW7unSnjugC
04wQ9OnEXPBkdGPK5v2r6tFv8AhJIEb7Key8vRAmAZg6Q57MTMCMjQl+YPVDlm5KyFv8r1hbc2qE
xIJOJOml84Yx9ZndyX9zsJ1+UyNNnAJ/NevVl7DsAiBBnBErQw/0ZnJID9EUXtvaKWKiVlN4KK+H
Fl1uuOYvzPbCS7NDg5MMsZqMBSAbH9CC4hi8YOM2uToGfPLdoRNPE6SmJmMAgvhWlcvG6UsD5pvJ
QZ/6c6f0T/dEZb0DxyUmNT39HzL4sdfdlmcK0cTrWzIWKtexy53coFYwMZ4pHC7/LoYkM9/EABJZ
VtojyYJ0k04rHhgeQCbla4lEomGx8lg8QF8O4o3uNB2ODO5OhVvtX1G/2lFDxPFNPZAvH4vPP8Uh
qSOAFJyOhJ8k9MCWBnA8DVDBiLcPu9Va52qA5CRoVgWxSXkjt39g9pDGi5e1ypqqKrjmx618YTkN
9zqj9g9p4ArrmOpn5EFtRQ3Gz8PwELqDBt3Gz6zUyR5iW+9dAPDyz7zRNMZ2kiyx6kx+XGAB2YHs
rsTSppPa5DpNHA2Z3DskG/ddk9xrvnvuGfXtUs+dgwpA6LViO8A9JjvW876p13m3adfG7uqB4m4u
SoRf/vwGYaHIE4BOGrHJBoeBXLwSk6kLdc+TSN9BJhDDNo5PTsmkaGDY99AjKxhlFkQiTiNOTYIB
nejTutbGCcporOTcs6IuO41licgWQ5YPaHRCheIdk/uaWWiQVx06kE/+HeyqIgzNu+sGbXnE/aK2
YRjTqOnkmPs0lAy8yYEBCXVbK8WzNXW/ZW0hM9MjdwJmx7mO400SgutwwPYH7/Ope5Z0Ag02LvAB
vfrFMNs/DlNAgB0ZeOh5h9a0elZIcA66acF6w9rwUK4E1y0zPsAUREF8kVQid6bPNQf7rIY37+ZT
yE918DMdMhmC2DTSO2LvU1siwNL8hZfQaPZ6d9d7wQdJnwmatM3Vs2GoIFb8zAL6KE+fLFe1zwqw
HegHGgMU/G4Uww+VjFRbd1HrAjy/+FLJ6ztHxMPgTgQQlqCWr+Vi2DA5+8keQcJBSUR7t8UqWVIY
siXhaVTEQ91UpkHXcQ0DPudLqkifMOxaLhQKOBaSeFmRPhFF8LX0XsGzz161i7QnsxpOLa4buJYB
HH1l+0cCx30U92OalEg7S2PhCkSR1lFMa2/AvJvpjQpVkOdAsc2CTTfatQg2OjGKWwABWCofLazd
5Zu90dEs96oBzVXlfeHzta2bWul5764rIwL6NQYc39VCJn2QV1XjyY2oddjeDlhJPy357/dIWX6s
ChXLfimRtJ80f9ehn17nsKLGMtIrEE53Xt4/MV3mKJdgktw5QXJL41YuQ3Kj3dZgT/MMeMsk/dP+
Ifnbx8T1/OOVgzw8MUzuAup7alRe+JpODdZJyfMJHtEVAwk9ea6RunkTmh2Zsab+X/ayBj8YJdAJ
CprgBmFzjLN/rO0dJ6X9IqD08q9w32qMM/tRgzhIUakYerC7mqo9ortQVOMGgrDf6IY846bdwBWv
Evc9F2jxD3b0eD1vxENyS8H/FB9p2xCS7Bg0VOEZ7GIA7rTfxLjzm17nd9C1EIqyNnKCn9MOZyUa
m5+kIIqCv+ALsOrAJBkWmJDLZgeDk2MWkBMOgAEM/G2XyVvDOiKcsfFbo1IoE/oMTDBuuW+vfVaP
O0nPljWP7TuC0ZqUXuRV4f5L6RMJr2z4jnuhKncNOzBdJuqX/sUwWfe/PnuOUbMlgff/Ka9vmhLs
DtcWliTjfj6XjP4nn8RaX0m1oM26msvEdfyX/ius/6tIUYcUT/PnC4dnvIfEfCdmLDbA+KntR4LA
pzaspoXGZgZV72IZ3DlVUF0wLoLPwTGfOwIOEGuoC8+xr/IouMUe0JdkfCyYP/+ojT3OrGqS5qrY
vQ4G9y/srl//el5InWpWEkUlV7nSBvp85EJxgd3cg+gxvZmwVsfh5xI9bhL+jU7PidSMXciMfC1g
R6c3NdZ+KGdk7c1rkl5x5eqwUMhgKV7SOk6z3HirP7wKbenn1sCfR/k9u9gQn90g6pUGdzoLTL2D
mRl2/sE2iO38MvY9xMqg+su6vwpol0wjQ1E+fCR/ht7B89Hn/6r8+kJxmpy5ayq/jZZ1u/dzFQo9
qieryYrvDH270J75wVXNrKTcwGZrAPQeFNKxY62v8gd+GCpX+hy+SJ4U29MsCPPjtnxK0MDfltCB
RzD+b2BHjEuvuYXFEhIf/9dD+tD+rT6zo2iyZRaJ501OuNzy9V6SrUfbTvKKJJzqtz4dcfGnydCu
EJDJQ90+YNNSbHx+2iULkhw5ctS5+sx/qXrgnWuwOCb/pPVHvDeCj9Rt1peB4QaS3Hfp2LgGCdqi
8RvsdphPV0Qgty8zQnlZySHl+IIhD+hLm6rZBW10zZ3J99KCi0GrAd1ufyV+lHRfNxWa9kDwkCfo
TJ3iCV2BwAd5OWHPQTuojH1GgSprxzcXh0kDYU3VZdqWMc3Es1NjX2qQZpF/2Fhm8NW64cLrzIc6
VKfRSd1G9yzfeYJaWTi4nWO7DiMBKcmKvQGeAX5j1kkcn6I31h8PlknB/F/Wd3fsNW7HUcvDSyx/
y7mOkXoK071SMVY6dokFwQKi3hZkZFJmURYKUUA++4YGpK/XQyMZEzyQJPXuDn1NaIB7bPmeVUyq
dz7KxqnFWpzwe8/3C6tZOMlU7szNAkE0vVtebH5VdRJ490mHwiDa2wZFWPYnCoh3bwus2hqlY+bX
QWvTuXmpjDO14UJegNyNMxtfHlJ52AsmLnVnUjs/tUWRiE7rorJ/HGd9mcurmdq/CrgYI+ruNGT6
QY0mz5rW6GFH7Qf3e3SEDGf0ZlUre6BZsol96fuZMvMRLWGzERX+wKgtIHlF7afAw91t98i3z/kn
xEScwrvdCq4+xc0r6xEeY3oCmpjm2qZdrlAzL1P5r+/YHBhMMScHi6EGninTlCSqOhumLpf6EddY
cxsIroRIF2Il0oDEFHhs8UeGS4UFlpDNIpGCcrztDrGTU5Ylj3o/ile98dT/OjzZiGAs3qj51Sud
oqy5rLBUo1o8IMVkmnIbysxT3VEDHki9npHbKNbIeCCVkk7YEA6o4vW3eO7EVyE9I8H29YDYUF+e
J6VwFD5fHUgB+DhTNeErbdN/EcS4Wtm1FqclwnQQMQlXlYb9ItKDDl5rivaMpKUvSCBd4gRglC7O
leoiiJhTmVuU+BA9H9/yLsb6zs5WgGZIfmF33kPmarSa39fi/oQuNZFnHV7Stg4KzL63HGSEBQAS
3RuONaIl9E2yS2kTFN/4mgr9EefH4Gfu4bjV1uFLILPzcoShESSGvg8+VkqnIWijA+9yGgtXzUAp
LhZT7G2rXlx811naI5iIPjDyGqSlBBF2aPcoowhhqsvXDsLhYnCzvBOL5EndFvcg7wSn1fuPtvwx
3zjerxaVtbKyHdtcX6MVIGvN3ETeCx/LM8H5GEqequ+JrObAb0QKssi5lZtsSLyJcIy2XPLZdNPp
rFEsz9JUsu12k1XaM+Bir5p5N+YHiqhNGWf9kulNaJr4GZDLBmBOJFrwIhN/l4B5wYqKGqfx+/io
rgpqwcGkVRw9f+cb5EeXuxhLQnWNB8AbuYeQuGCJP4FPxjD12AA7DaNrvEchF15JQMKuiAfrJsAc
x02MJsZhkv0XB/7XEOn0Ptu8iDcClHVoAg2/MdRxQ6a1Lh5E0UZ0lEgbIFX5FEvJnI4zRMuH9mc/
ovB91ARxmjbiU/FewjrlqY8W30+f5Hx2xMRhfcD1Ymzs3vcp55J3zQ3o8bPMdWWu3AYEkDapWlho
vMHu+6oyfHn+v/tV/uGcp3tNKRFTUhz2U7VpBA4IgVJMkm7s9bRbrWMV0SjK5N8SxqAyU5JaR7hr
RLmOCuFGduAtJc3OMcAkk/eK48v8d8/Zk1Yk+5Vujdu79zNycp53XrL1Ja91kFdeoQqFTbHtrR/n
5ueQjywyBVdo9HRAQLZeG3shEt+Pf/6CAnwwx36W9C6mw8o1x5AdniBIH5PeE8qbGtlvfj6+DyY2
Mu+Nx43NoKdeUq8fdvrAo5VhEYdijOFul/0CkMiHECCJVAo3+R9YZihVqrn9Xu1ueQClUci7Ntoh
GOOcG2QG0YYqjxTOeuEtlNFuuoTG7SvqnH+PlGm2bcMz2E59SNxlbm8gMjRHECsjozpBdzA0geOA
DWynwDAXe6tioLEd5fHEU2Ps7neOlKvODQVLwBbO3BpZJpLv0t+jGuphOCfD0lsvwaEYL7qMCSEM
CI43mWJ7/AtD8j6DEKeYcT99UAP9q/6xWoFz8GGFeCHdmhSHIrxL//6EBVwg3yjGPOoxiCE0dhoC
4yaJ4GzZgRvyQfunMjZSntS/WRbtceWKbRLcafObbov3QmBYgeWDS//Lzwn02o+A82tjlWW9OOQR
rVqWohffGqKx+KqIquaHCZcM0n22cdPeCGeihxBXLNZ7b5u7jBP2IXciFKxgDxvfxislnrGB92hZ
h3Eu3YUYVvG/U0dnpB15DuP4QFdcD9jCZ8eLubqGoMh6F/0bztkD8XDjPXxn5zBvR0M4vwp91bXP
5FA2KOHQskBeVrfWX6QLONvUrTt/7lwS9srVYsgYBNaN+DmLvKW5pg/gE+UNR07Cq+kU8cgEt0qZ
ByVRGfTXv9Ve7XYDKrzLQnnyBdZVSD1TiffTcNzmpCjg6s3sBwwfSyMsmj6eiiJj2KPFR0tGY2Ro
hPCkpSqV0CeeoWKeBNmEzzz0JJJJ/Hfhuvbcvz+8w38+foC++OxuHTij8l9xYb2kNDDjvJBz3Z/R
WcKiydIKNJKzNsso6VarBVkUW97s9UxLClgwBdEDkQMiG3Gx4oMrCR9hCiEGd1AmFbR/RpJehM5n
9ZH/56jTKxjH2q53+6ry7soTzZz53zcBSUjyzr857uw2u7MLpmc/vUkEmZ8v3PEHPYgM3S/tarXI
ejlL8XGjJe2jehFKdOxNkbllSRUEGs/dcPMbTmlvkcylsMCnHdgQPOYGMbLS1DERNtmw3S4ToINh
NkZzd31x9TC6jf0JrERauNvH6ZrviOaZl1HWtJcvIbQAgBL88/kDLY2Osn9zJcBAADByMLzvofT6
IAm2ETLf5SHVpqs4mv9k4nXaxjo/j74aGtq0MahXtwQ+aW0hwFB+0L4TyFHjFCS4FvAJ9U3mldgh
Yx0r+6Uh9WhuWt/m2G5x2O93ogxVnBhEVrFf4Cn3rU3fQ9P+fppqKNsha+gAXmn0pIxAhDUNQhN3
KfqKWX1SPy1sPygrFbNAo3dVDqBUbzPVDxBBWfsKLhFwvb9ObuzOTLWvsyV+riFT2jo+YG5t97fx
D5iAGBzHuI0G+ZW6qN1p+o9aFt+d9501gfvpIKJTpNWZoL25D5ff2zMmKHWy30O1TEf++dvmfu/I
EoY8qgyc96+N2wzIbmU66rrGB8F6jdRS37CkmIyu6X0nyoDdgkMdV/9h5haFiptYR6KKuU0EDbZO
xdVPNQI/b65M5f76p4bTYJIHBwEoCTPSPoSzi3SylsKqaVRhjFdgRiFRoN7Xn8AAW+iWY1IYeHZ1
3ZGZYV0KRCFlSHyVQvMvfJcOEqtVBGfKCdNo9TDeMJn05CmSJcySU4XvDbRGVAqCsUK3eDkdDNhO
VJ/b8FYSZAddDaxjNtQ4+v/u1NaIPebl5cKyEifs7FETtmKtb8WGvevZtmBePt4qfeUXZ2ybJac7
l7kh7lP+88swlQbx8Cuc4x3VgHLOpdUk6BJ251+Q89Ojh1F3s3HK5xES3zNOOdq0Pxx/MuIbTl4p
6KfMPiKDjNu+wppOtPjKoQtYY+BAMne3R59nYyo17TkkL4FSCfu4byO41d46RP94jA+Ij2nBgoNL
6wK2h0s2THe/xL4tbPkqXoSI0CpkT4fm0gRhTatZvtGaS4/R0v7TOFD/C7/Cf9euD9wDjb87hxhI
BM02OJZU0XAEkmyH+6e/w/S64BnqMFh9pPFeuhFgevXAUJJpGAKBRX8snfa4Rt+fSj7RgcMM6FDZ
7awvgHH5Ik7Fn2KZx9nmznlsKKg4XfiZpZolDTwGIDWhkYUbx5v9U7F813nLWhmJPfqe7HlHmSqo
Kr88PUTBzSD7EtmDaPL+CQfGqSDjda2epcV8wmyfx7j9J4ZNAzHAbl0sEIF2w4FZuHytpfuNr52L
vqi+mUgrNZhLCeXWtKavhJToeLSfhLJRPSt5Iex4PzKIi23X3IYNb5dA/ZkYHu4Y2Gr7UCotOW4i
gckRnTlZ8p5+JmjdRDEs4ojcPDa1k0UR5fEb9qyir6QedPbbT6M4POV78P8iPvUlDEOWs2LbDmEh
gBWjrr8PBzFZXK4/3LZAV+JAoc4lW4MkjeMHujQ1UisQR0ZZ7Fxj5fhO5FukxzsqbBMMJw0edU88
Bh2FRZ2RaRzn8XqTwq4xZPHiar8SpkEWDz73T3BJqcJJ6lyHx/SCxWQ7zhah8HFeMiaw09FSsASi
Ume4/gVSz2Sz0lxGIIL4ZmIkCK68SnyQgyciO0pfGk7N+mO7x0UhsFr80BNh+Hwr+Ow/strDC567
UgIOGPpBiawAdikhfiiQIapiSZgDVX1Qxo79HdI9VBfjCgpDTJKgCgzPwWpKdpA3szaf63b7Fp+S
VCMo6cjkp37/5oRe6ux05iWfBiSG0LVl/RHAxiczZk/9t/tK0giiionhjT8P/jy6jWOo0R4RHKjm
T9bjXJb4OfN0CLYlkTjgF70/p+CJVmx6Ep+EvYYTvxP70lL8hsVUWB/eycQ7dQ0BAj/z7PjHZyW/
6Ee7xukfleiw+CusYLVW7/kGRR15llzXkeIqgCkHSRSJCuF+gWt1LzQYx0KtGIcauBZMd46zfERB
JYRwOJcEvpe1WZhPdkQus3AgUiTDgQDPOSvqlQd5dCfx7RIyjeRpJFL4ao1a9zBbgUduiLdRbBAJ
XDpMZFp5v23INw9xZoqloWkS1B61u6OmAptGn1zlC0YGvzDJi2OhyxosRdoOQDzzNcXLRv4DS99f
FpDBojX5ybx5ml7g71vmTg8ywY9WqJVs05OBohNYgti3wIbsdPcuiPmrdBMFcnvsLYRsgMjn/ErW
MHcHHY0UuBRhEOhR5sp3K1uI1iASFIniHDqVO5/Xn153SELw8dsVjHNQPbSpDEY3Q8jQUxNsmRyF
vtNGXCY3BSUCn5tx9wh/uAOVld00NXKmsLfZZ2QwbDdV1ljfKsmA1D+emnucdhPTPNVzyi1+vVVP
VVWRfzrNvT+Pb52G47yQYBUjsOkd1tQLzhE1yLGvAfv+opVN1Fo4i5DP/KoYNdodl05F3P28icyz
myKDI0d8wDawPzOK/iHVxlCBTKpOGHE7F8Dx/OjCTUc7I3YjauHFyTzzhPtjABR8Aku+3f1QBTnq
HpNqdU7QhseC+zIPZc0WwnUPcpYV8fGCrKaLwd9COHdtbUE8pXaqekPMnYSuB+XwyOg/eChS0TDJ
v9dUC3T5IS/LwDgo+PloRrjN+pvh4IJKTsFWqmyMLWkwSt9ubPuGeMdPSG+AK0vhxEGYaTyIEsqA
VIP+VplMotHboggmtEDAGlD357cLpSrgGBopK8B7HQVvRa3MRun98r/WwyVvCaEM925cM+zn+1ET
hRNU8xbffchzf2MUObcZZ/skUHpxecKMcVljsPc5ZyrAPdjMp/dUfwANRqaCjo7nJWJYIT0R538g
+QftIQ1OoJutiQMGvEULmkT2ayyAKr3u5oPeX7S443LYXN8jqVU68BU05ATLbY3ATR7nRc3Aau17
Qf5t47X7M+CgX5xK80OYsRKPXdWrkPmgA8nKzXak6djFr79jUZaNeIfFIXWLWSM3iVz4eYx/ouaY
bUUhP1JWbWMu5oFxutjAY7OI+XO13M8v+5bsvN7XyA17C7sjsWqyK5l3M15Q0Uto7M17vHiOd20l
MskjljUMyhzAPuBFjJsSbiwqPS9xyT5LEGr0thESLmeljFtxGX4AvGjRBCu8kPEZygbICXsgx/7m
tNiINKUkwGxzKI1kri4oV22TG/av7HeNz0cNbbRcLDnm1C3LbyZHjfSkO6m15akcRTHXHU3gR90g
+Bmmv3a96Np0KAzPGfskNnuQMxD5/sTQB1IrUVJ8D63WTiZZXrAvPhLyHpj+RcZy22c1OfHfG424
LNEurId/pMNAWmm5YIVgNx3p+RjA/K3Fa8AuJiFnEt41pzU2bENoD8iWMfA9pxaT4CSrOkt6aCgN
XZbhRjXmcR1YuH+oVUYmPze00yrkGPYHjNVww8vryX2ZDE70iHV6BHtAUCVLIfw1j5bzSglL1ypc
JYWhdxx6NpuFC4CZdbsXFUHlvjNKdabfgfYjpFLl4Y4ersr5tsr3QBgMezALqLcQw3HZgpZhPPUe
pLLMmWuD1YswJ31MXVxqywcUoocnag3mRNAgo7wJdQ+pA4We+s9kUO95GEhZiRaObbE6wCaNPhHJ
3Mdpu4q51BMWY6Xlzm6vY+mgvGwQvdUMghN+2dQJA0Do4iNq/Bcd3qdgT8S/9gcRx4/L7Uh+cnaw
QuPoXlE8IjnVw5j3WOcbglKfyhgHOjYrfZmJAvHnKrUAPhGxQRqeT4+NXEZhc0LjrXA4kEojpcYB
dxarRcpvf2Rkoyts4MlplEtEmI6sYU5/mmhpAAHhQcdyxIBTOXKYNYDc6SbUkoj0tP9dV8Rp0/fr
ZGfHwxBAVlyCmMRdo25RpLOpP2ezGXNMCG8pxsneJDpHZc9Sqc1f09JMbUQB6485usmU1Ma7OEsy
6uYSpOBJBbM0o+7Y+QoMGLJWAN/p4RL4mP5hHzSQQd50AqpnjfiBrIbMZeDm2kBerFtxnH5nNpns
XnSzO54NGYRdX4pDT0OQYWkFj5Novr1wtBa5KLq0vqfB9azxENIwFj5qu7M8CK+33IFzvzNLeh1d
1S47q+rdfs0yJ84VmR3GmCli7xLJgnXwD06wXZhohG6Q5kiJsC1quEDnsH03eIybDVjyn1Jr7n8y
d1JO8Ebvdu5MJ3qKJt6kYN84tw/fc6GKi1/gYfidA0c5bJEMJp2g6KgiCgKW2BSecEI+rkdmb7w2
ShZILIKU8alBoScaxEAAhQFxEC2nxEZkp7jNb3W5Gwm7lpfyw9MhgIl6yjFDz3J+mPOvSU4cO0DU
RKqRPMgB+8XKCxt1QWa5vAUEIbcvClcYjRyNAxQUCkpeBgHDOKULIZR3vGxyA6qPWEjjOynOhdHY
nZTO5CHYIgg8mFnbZ9/orqsiNLEJY2r4aPSrkxvUq1o1ODYKQLs9LKrbAH8IfTSgu0XSSflEjXoL
sb5zc0S3p83vZAWtKe6cTAi3041sf+rHksphLaKSwyjn00iK0mQsN/9e9V8iYFFToECMYXmnV4zk
BAgQXt36rnAOzcXsYR7ZMKKeFKam4vMJMgiBJob32bJfGDO2lwjDLcVxopozTgrnnUr3wnHcBPvJ
JoSklPUH7m1Isbyoxf3ij7/MDciVk9GiR41/gcLBPNJ9VjJ/rbb33peJAkDcdy0BCaZzecdIHwvh
XWrf5xx+5j9Hcgir4AnKPukMCVUAxj07XbobMajDWbAxorUdn0eZfRXa0SAwtkXyk3vGmXLYqfeF
kzToAdh1K4nES3+A5AY3I1aoq6ok1JBWzQy029EyRxmfAaBbkufUFqa0a9pAXjn6duYdVvg2Vmgo
5l667UjDQdJZuqzBNr/q+an85oSGWLKiVRHsatv8QENBk4xsUs6ayScl7Pj0HYA/iaEwtLDkXoF+
IZQQRMLAf82Cp8cLvO2oRqECMGB2oc8sFw4VsBccynKcN3zhlxmOV9hWDNMkGptFP8BIBJXOZd8q
Rmy1DQAjbCI+Q75s5UmQdamsG61u4dJFW9ItgzIMkH5ksR4XlYCSpirFCgdRwOwQ/PjGkRLMdJKW
g/Lv0+HWOYwFvNO585T5UvvQHGAIecBLV1RvFpfQInpdi7tN8qMrfxOMB+kK8zyYiBb4tJ62MT5Q
kgcQDpkN5VPh+OkaH4WQvhkXXdQKZp6+oK1QZgBDkn9ctdMKwdYToBR8VM2oA8ZwtZG1r+ivhggS
g25nn2lqyyNExQNZByjF2OBNrJtkWeCdG4Q24pz/571pDRJwyRimpGMDdSC84BB1/Prqt0wzx+JR
HX9+N1fPpejkZyk6M7+mW0b3QKkKto+EgSYKqJ72hdWmg81mecj1KNKj7usI3FWX/6neWCtb6gp5
TvfaqooEJ2Yf/UD1RSHXbVZC9MDht/qf7KCWrz/MIxWOJE6iaeLUPJwrEJwb8c/tSNsjl4AU85c/
o5wFdhlyVvX6hniqUMMNLvXlEqM3gAP4eQyoNUm85u5+ad3QxhjtlkTO71PXQydqg6aLH9qosVL9
RXEwQ5mokgOB3dGfKYlsjL1KtSrp9+Y+BX5T9N6xXQqumV5joYY90NE+Sh44giI2CJyLTGHKsD+s
uld+A3tq619DneQRn2aW4pJ3sqqS0D0DNq4AzWJyahbchCBBRb325G4SD/kkAZvB/BfAnG2hXKI+
tgZz/ZYhQuQKUk8/6egktynZe0mdQfHxhmb/ojAjY6ESJq0IU9YBYuo13T0bmzM3gyg407GLuE2g
ZdL4axnFblDrOyjlMJTCrBHiojS8+Yyy1Z7mbWmMPhOc6SWX4Vb9DVul9bAzLk+/Avga02/5Io+k
nvnEtbfLjZy7nHuozU7McDdgmj9fl/YhCIGzXw3Y6RJVOEogdv7wMmidIYdjgKPYaVHy0urBty2g
ESe9gl3W4kkaJSaU4h7IAwtpSifjf/WTGvqXhKanCQa5ucCSlma+Z22hJSNzADL3w07P8wLuJKbT
LdhOYm93WJ7HPzAd+XwaT8P+msBaYFi6vlwRfcnz824rpAi0dL1GXOdf5vXiCzt2affcn9JCJAIr
Lp8WwyyN0WRZVSp7s0YDY5MkSKupSkqlbwHUfvvSAR+iAPnsNle+yaDfnm9SO56FADLnUOqHd4u+
NGqlbBjAfnT/6PDRPBUghQDI43DBj2MzkFyDrDLuypeKQq+EAz7Syj+mLn5Fr8VHQM5eXgTta5IR
TBbtFNYeD8bVMi+Dvt8lc9AS1h0040Rjs/JnzC0eEQVVmxjktoSGRpZ2lLCirdJ3miyKvBPb92Ij
2iL2hofSmRebs8stdrQUyA6ewqwiC40kIl7JY7Gw2b/FO60hfnymaK/5vFfY7iRvkRHnOG64bxcC
9ZYvr4LAp+yeTwEKJf6plT+VRTSiofRFwxy3BGa/Yn5IZ5Hdu7u+ShX0qeXqfK0dygKYycvUG3iM
do+UKhAPZFRElswuz3XOS96B939Nthqt28WOyG3PbEB5PH7im7ocZ3QW6tcp/RACttBk5HO3EfVH
pytrfue3YdcvSUDxbwwWuOR+d+GGisBC8/YGIJTzQaJzWIzziSWzFbV8AIRanws3dZTK0jDs477j
Ctg5puy2e1H+RnCGzWyT0fQ+8CrZkENspBSiCmeJbhk603N815cG5CR4Ak93pwxLhtttwKx+BdfU
Cw+YpvvnYNYIEvCkB6bMO7LKZuO9aHNrAh2+jr0qd6SSedM/OGY8IvJ4ap3VOeZAIR8Hbara6pTX
+yM7xkS9N2V1iazwTJjis5RRx68UdQkeYyRn6YA35wTy8jn8t59tlGmmMOEVoFiAS3OtCz5ezkvT
FRK/PdrfkPQ0Z0jrWdxPbfy2xTyXcndJcBKTWV3gPAx9WnEBzwQpEp5XPxlk3/CICFL1lSGg1dSf
8ihIvMeHIhWA76RElJBlbHPMmv49qQE4AOkz06fn9/suribbtk2Nq+8uumpNIweF182PhxGzjJbL
izOa3fpzQ10U710QB69ljFXVfCrjTnZG38xbMW0cRGLhEtsuhbITAJfH3RMNM/rk318+RBksS4Cj
94lPMZxW7J32ZFTv0cmz2zW81VyyryWwzvJDVPb3KTon8wgStCaajo6DUWAp4s01cBkE2fkJfQ6R
B64sbVf/qJHG2FM4p6cADt4BwM1bB90bFBTlZ/A75awU8e2PNc2XohWEMwrUHpiFMq+gamVTQXgm
XY6kOvBUxUDXnf0iVD9lLvm01gnmozSZuxmqfLhDTvgnHq9voHZqGM+TW3qDgcEfCH+TetXQCoMM
dwuPRKOl/NKyCwfjkflBvr9FG4zMt0b3POJCKkPUe0mpRbryBHROZRNqQrJYl9uvpf4igeZlKlZL
XovHcn7FHQPLBauSpUdUQ5mwHMye0rUGI3HySAsOzitH0UpG78J5g2dkVLxQsXoTetcQyAf7eaZC
EnuN3ReagR9OJKCwtH88DHWkCfPMj604ByhGXe+A+df4I4d3ZoUnkLtF2RhPpyp+/Ax3yHW5nkUk
ieXvi9u2rzIkV/eVKGeX0K5Y2IG/C4VEhUlEa7vcOruNA/tPseTiGup0x6qYQi2WMz33N17aCAko
iwJWu7KpEUFvRZe6KWDW4erQnRCW+IPEijRZjMB6zILNQBDHMdePbE2uuzLg6RAVBvv9FtL+SvD2
lW+TF8nVx/64gHr02j3pt/j04f4f5XG12VMj52J/QOVBQQTEhK/XfP+py5Cer7w2y7a1m5tG1IcO
WFmSH9Vs8QjP4t56LOCjOsiIarYtLWrgSW21OeN48vdUXOthy+t6FJcdU5bCBP8KGNFu3e1/uwtF
79FjxHOtG0bEEAWpLUJsLS2XstvSIBeSfXSJkI954gci9ispWpOKzrVYMmdGRrQ8x2o5y5r7sGPT
CGiEOeokIJDPJIAguUJOiKeJLnIxMKyk1R9+HI4E8vG/jFEEMHDp91CWcPMjIWXFMXAXuuCg0kxt
aOInxlkeIHyDW4+Kem0TaTz/l2SU34UO/3f1ZObvfj0QtWi4WYUAoaOFXQngtWqtUwi7YnthCvjx
lH0MBzKwfnMdJBcGvQR1wMA62JYd2HsBIofH4UGXusPLkLZ41dp9zEZJDxbknc8Iw24+gzowIg57
i808SC1Be/QuwBPqHXb8Tg6A3rO2j7nA/nPjlkfMXruWIQyZtsuFdYQ1WmAQsnUZiZlnX/kkMwia
Nl/NuyOTOk/eCpQh+OLJ7J7wJ1fXBMsSEQJuh1cKcipox7cVwW1Urs61I6JK0exRd7/8nT4++KVp
64II4B8EZGUHW+ICazBWrILKLN57Brg5E1OqCZM+tsdTIlZGg94zeZDUZfiv3NBGpf+UOU6tcIst
h7I4adFG+mEPBJA9TAWvPGnTtjh9+v1OfqqANlvGMYIFn0IHoLEWo/rY8w6Wn0yCF05sSjSrBqJ4
+hUFk93c26EawsQ+9U30ilEf5rr+8Fz2A4EgJZ8g92mMUbIdG8HfceR7LN20lS0H7durajpIuQ1M
uagZg33O4Eao56cNRP9qNv57LfbPa7LTp9r0AXZwcwwvr/loNPH7pgejLQcQ4rf+1IJsdhgNYgkP
1u+9nHbLBrWzKa9irnbdMc6CcxgC12sVBLUrICwb8cZHrlPc8o+pO0ejrao261yWrNQRzEbKjy3K
qC+VE/pPH8YceKNOPmDRr8lcR2uVxSGxryTSoUS3orb7aAnJMuGnPf34i36a0Czv1txFaYASHrrS
Ou/96RbcCcCF++Vne2xdfKckjLdYHp1MZ32Dp6JTdgGq/uifJg9ik4WiYN+qQtSa/rVhQhh4KVZO
fPE/aUAqG/ROfJmI3J6hs5N5FD2ns2/Kq7bHr3Pg1tq16Ddx3gUFhRsqdH+QyoGjiAb072u/eVWX
15WcsVf6ZZfbgBxxmW2ZxRyYt+A0EqeMHpJT04hNLZsrT1W/+6xSqFBAxNeB+uR5YwnT/aUS+yB1
PueOGMZdR8RLQNWPg59nxIc7GGuGJC50F/nr62knzt3Wm21y5cQb9YZDg7XxFGXsUIo7wxMzebEC
l9Kbgh+sCKG9ajqB3xkXHIfqtNDOEK2kJULwdg2R46utonN+dURO3ruXPewIjdu9+6VJx6kJIB+F
hFkjBaBdhii62A3Bu80kYUbdl2SKopqp7VpVP77+hokwOIWLV5ijDbA4FCyXxGoU59AnrogBp7NP
PXs9/qWUXQtwbisYffTRmHvh4oHcDVe+2pSCcVWd51lMFPP/ER+o36Z4DqBaWJsVgHsyfJAZfhcN
USXEO+9owSXpJ3H5cQCr3VCgrhbYW9zL0nFz7cRTKTZeepqKNJt2Hllceq8LmxfXiXQE8dl6sivk
PQVlWSHAaOw5zQ55df+/lrhjiyGkySt71eheLoKixecZLraow4eDqQlqyhYaPomDow6FZO2myVfr
WPxWJsfl5/YTfBtcqwYodFD+9djphblFmL6S5fRT928qotyuOYy7RTEFcq4+a2NPNFfnZkiOTfOD
YsytbI3NLIxLkRJYDVqQeyapItffENmjhGCqp/tjfCUkE6fKjVG4eigEt5/jeTLffAmROwGsw6dZ
9b8YuCwYnJpPORjhaoNebnUnv/7hGL2WkHpCheZ582mN5zeOiAXsGTCVBNMyfEReQ/IzjmysiA7w
jO1njfu5NRB4MGDfzOJUyrn/WaGqACzLJ7RQ4gj58d1gtiYasQeQj5/kk226prNvmFHfAxPGH+jt
P7WNi038ULjAXc7QIFOWAd6nM0/qvqEvWU+aPsA2I6NB133tIhGgSqZjBm8IHQIDNCkK/I+NmWxp
aX7RNJRJwicJZ9wUV3R7wxE6B6awmmuoWd8v+9Ug/uAjXJkENhJDxDrC9BuULuoOT8283VSTyIPi
Pcjci/f0Z9sgTFAwLsyxZh08V05qV/6yodCbu03mBSXq7gytVRcyvgG/KLbOBJ9oZRShHXa22HxY
vokdcYIXfTiQcVVJzdGMYq532X/gGA8wvrys3q/jdvZUNSotFKCSlg2dz/PzGMQcs9xwODefky5/
IrAQdGZ4nz1HSkaFuJgRHeG4/KCY/pIZOwAJWk9216h1UXEHdjiLK3u3DBBEdE0WwPdsci9Gl9G1
qE0skwVSsH4ymD5RSlbLgKaXyG4jDp96Fd9vG4e+jS+rad/pmv3Q/TxSAbbo28yMwIHtGdwMSDQX
QupsiQKcVnTHw/b48AxB38u4ZxzHTSSa0HWm2JYHOyZw/z1+qhhsyO38Z/vTqiO4WLZlvJESNeEs
LP9YlDIf1Tqfcr+9p80c6mjkGpfJeuCnJx/KewHJQ0PfkNttjWd4DjYz8ykwsQoeYknPtflRjLq4
ZlFKmHDN9Hg0axxrc48nO9QiNMgCzYBMsjPx0anmKOsoV0tQUqXSvsx/qW4MJZngVbhRkd+hZs3e
Im2e7bEMPF4d+fJhgc4rWm0lQvodPb2qweTiN8U8XUReQ1//Zcdu4sg9pzFFRaYHCkfxQlw9Tgey
5hPmmsujwmT2YQIOzQzlJxGnyp+0+/KYBHI06AeaCYviS5ObthZ98iIRn+svut7SMjsqtJwqQ6RB
rnryeumam5Xih0XEIKLaYN596LrvUDs2jlLbv6R3MkLM8PrwvLd3OYURmW4jrrmVxwj3kV3Nghlz
bnihbDGoxZXi5Yu3ssbec7FPxPhvWBbjVLpNqlA7hmf3TKEC5dVmvoQL//G9iK22vSD31INM/LMR
PUyQxi6KTgP465EvaABMnybOQYBV+thJVGRRBtyIyXNZo+Zi6DWaiRCVusKcv4zeJ3Vw8joRi7EP
W9mO4fcLIMvC4glj4TuL4ErNsbMvmryR0YnNZdu3sxMALA/6brDjXwXIGund02a2cGiOw/y1MusS
XRi50frXcfkuKoGXqgxiVgEkhTZtwnLx8y34d9NuBNSmkM/QIkEpmJv52xqUNLjzWwpO+R2emnAS
Sk/gGOsQ32eQVUOsxdTbXZuysolH9PksVgpy97ey506H9lAiSDRCAahABm0VnQorIrSZsASWoZeY
HGAROnB9OGX3+fKvWgp89zOMDdbvWJv+0xtuNTKVMrN0kKoZuhgMEnaEQvw0tlZRCa0171sPdPTJ
N9P7lYSRW6VB31Vm/mM8/LUXlwtYQSuA9d5m41ipM5FGco8+zQ8SLqQfyGOuEkC3n0ehqaOfZ+h4
ighr7lHmI+felfl3qUdTj8aIiPGiU71lfGKaIg72n6nzC4h+uWiemnyZ04SF/TPWwVkxoJ0NSklK
sivOD972n3r+3sn4Azb3k3Oz4EwqamGYjCc23LqWt9szngrJc5R1I9+H9Fkpe6wNq4p3HIkgd0vB
kNaBxYC12cBRB5ytSjuKMczYIXWB7zzWM2YsT4yruyW1qUS31Rrly7a9CoNnoHt66o5o8BjFR6/I
Mix0FwjT7mAEZ/HOjqmo4PeuaZmb8q1GDYiD/rvHpnQHWRCaRNFyIJBj8qqy49uXwHAd/Pe8JYwq
86hrqBEBykV1/N6LENdsJZZH5n1gUZHYSaRgzlin7PupxH01wazQ6tagu7AlSPk8gyqzh6RGHtYs
S3eg7WRAQYr+InAS6qH15SNdQfw/u9kmOX9CWC08XNf0ps56d/Kg8Fh3mZHtQsCgKPwvMr4m7ziA
t6a59Xq3CCHeLQ3KuqHYgWQyHhwZBx2O6dgPtA97FXCpsxvG4pdTiu4kQz52ZukAhKNPPSIdD3tH
XTa5K9+hr+iNymA8YILnj1mvkw9zVMeQjvYguLKkm2ozoYhuzwIyYziI2a/McGHMLctXwv8HJHkK
7wENsuXLoh/X2XyP1X3ABtSVfn4MJCUFoQM7DuTAmPpDeiB47PG8SoBkDIvN8AheA/LZ2DGTzsi9
xL4uMQ4Ysq1rHSVUxEBhPeH8sonvW+ggCHK1205r130vRLqGbKgvfDa0o1aoF9a2ni63ddzOBSnX
KgNqaNkq+z8wJr2E2VL/VEyINBJL5nWZFFRu6WHHhTqbEhcDKLbDBA4Fnq4QnnGpk9AjifFV5yfd
B1MRSkUj9nRlYBpCKU+pls/sQkKImPaOzc2uKbBVQUh+xM/KPK31ym5vzqc3pVTzO3KF4EiXX258
Qxz+4YGI6V4DHWAA3uqItyUZ2F5Ia9WRnrSW2oRpD2++ME7ND9aL6hbs5lwbt/NE6bRM0fpe56zF
tyGFrSnYmSXxGJAMgmCEaQCXWOlmvC1mRGnu30oICIzA9fBmZlON0SvP4GWUv/4SYDiAI6jpflFW
q+2CMwpVJOjL0EezLiDFIdVZfS9kl4QGPvTxQOxV85+HOb5Zn4bJR1jKlnW7Z4mnUmr7EZy/mrsf
vjLlZxrAsOGpNqJgtdtC70uvl54dLLqKqlzQKeIKMJ4gxalR2RmhS7bZbaO7H1TiPrtox0ne4dQg
pW24qfEkF2CheAmXyAOIRe2b5ebn/Ae9cHXqxZVh7Pw9rY7HQ2aSwiiBiaJ9VY4fYJc0RJb1WJgO
vYbZxQMMD3gHXTTMq4lLN5IbVmFetv2zM7U/aECRRIqbtygmg3vOrh476V3fSERKYD0GlM/L1n7Z
V19VT8mHUCfAmbhqFcucDWol7KbNqw6Qa+Aw/EFNeVD8buRopVr8ZqTj3NcD06MOHOPj1BxLOBBZ
ap5qpWv4LMREHwVCNwclInktJzFss0TEymKxL5jzgY5uvMSToEROCzMY4/QftYvOXkUi4/xna1wz
u2nSClwbpe1JMsN89iOSBjgcBzX3xuuqAtm2ka14Jl51w9nZ6JHomglhzqD0kF7NDe/AReElK8gm
Rg96y+dRm0AsLFk96Mxw97P8Fm37mQoCpfoK005P7UGqS7W7WH+kkJa+mw6mqE2pzQzAQtZ33TrR
iTMSC4KE3It6egeYePKXcrr0wMZ4gO6HCwIlp/rZJseAAHT4fd0jgalo/ygGG6sxtFIdqBufrHLM
g0xoaLYM0nXC4WZKF5RF55xAcffBi+iAeP8kt3XdNwbZZ6Er5nJ4yChbaoLdQERZ57NjpPfV5ZR7
OzU0Gqk4J/B37yfx0vOtdCgJnqdIdY5Ti0o4+QCKmdBPtkI/BqoRRoX9Y/TZWGAe8JCutz6n/ra8
512ZP6Sfre7oR0qQtHUkr/Zn6MWHdnfaavJsp7hrqjCDUAbA6Z1qX1FD6GvKrpzSdAcbyyiC+9X9
TRrM5gB4q+WJ20pw+XbhmckscShmiAGs4yhiH0bvjPrBXzZ8i/mG9vyDYhdeq8Ab1x7OzqgmGPJ1
+HIGt3CpF4aNImdG+8cR1eb3wSyT1v5x7l9yEMtn4IFNL1wr8Fbsd2ALhvs3ioexS9yxHhFBSURf
+p0ok+ibc7T9mA8UvESk9OXX/bOjxMtq2l0cLdLEWKq3BfseFCWiXv8XHLvIEpPVZGGPF/rvg9Pv
M0nu92vQcc1Zf6cR+Fum7htDFloglWIsNVDEYvf0xaf13gEseJexyJZ53UYSw5rRATa3P+3/dqnQ
6X8aPGhJZlr5OtCqZIR2EX1Rt4EEY7TNIBOAhlcbx8ZwX6W8QGcZsdytpY6gFhfGd+L9MSCbF/S4
A6M71nUYpQTgvNSCYriS8ejVVUb5lvYTfU1OQqk4c3jDACj+JaPULqTP4L0MfYoJmR0ekNdSCg3T
RZ7zXDob0Grd6B6HagMuIf8xdk8rIdoB2LV6Nbvl/BAuplk3hAZx/UMFWc2em2wK9tdULcc8shOO
Y2F0LfADnUi/mvNSRRNfEx59oADtLOGi4PuPp9uWtNN1n/n7/4J1VWzSRUS6uqX3bP+Dy6z8Ve63
4hxJqpq/gBgd9qjznQqXqGv1uj4M0g80dng5QGC9zJtFiSPl2CHZVNiBj81PGPZQE31O8xBhSQ9B
JhhzddpH5WNpEkzpweZM6X6fks+tKauPz281lIAPK9uwN8k1zM19QJP6i8hNV7Uyt996xc7zAtal
KeUnU8hNMCKn4vMqWO33BzqW2JXLtwe82Sxvq0oUQNIHwSj37nYmpZB/+6AzRr1J0C8SfXPL4TbY
mtaGfKbv+RXkAlOCqNV5czybry1EM3kGeXhnYCxEy0WIm0CHEL6Tjby1yCVyhGsiQUpZYDc1RaHQ
rwJxRtZGW3l5FghYc7ceJiB1/yeKSPUJrR+PbqHTXac0AVniIY/GaTrhgkV7n/di+E7tOoskMoPY
GBx74epwoGyGHfIF1Ul2fKme3nmZMsJ0wQefo9ksWUuHn8L7Ww6MlCctqRhj3H6/4ZQJvayAG+fz
LCmFD+ffbOqWhkW00e7Kdz8oMEfku0Ye3XSnRfBr/NLlPiZkADeyy90TiEjDNmsmozOb1IZXazFt
T8z9PdFdOo9FomXTyw/s+khYZOWvRuoV5ytijxkJvVW9M/CoK8Saw/LRABRZQfe4UUacHH+/4F4U
TlFfDlNicIBTh70wOeOnlyxy7WEdBGNeZsA3vWPXYuC2wgxC6g4O1XnyD41WPp0NdFFrb9JCGpOv
G7wH7WR70UbcWRNFLO2Pg1Ol0Zmr3hTNOvjZtfsEoAG2yetDU1d+2agG5NT2cxLs7KFYuJaT7cfw
Zzg0p5I5/t7UCH/KciuDnw/jB7R1F9W3Fd4QlS/XpXVGZqP6Bnt5Lg3v77YLn0hMQGKO7dCWoF/n
2//oXeDaLV3OZdFDvQS/5n4zBnuEA5wB9LjsE8K5hT8L4xTwSwRvBpgIO339DI1wf9OBmfvmvwOC
UCRS9AYM0CS4wkAPPZc8k2f7ixHLK8yGy0rmKw1TpTMRTHSAcmvogGp+2Wx/8SDl4uuVHaUPUqw3
IVMSdya75wr//Cd6ulFbTwDCpbtqhg+ZOHpRZH0UVqK97BGp13e21aaU++4/pDmeAL3itHpo6AGd
0WR1R0YxIF/kkW2PP0SAYCF4Nwmf16TGqK+dXgBBofb9zdH1cs24+97FdPDopKYsPrWS2IAZlFW9
XqxPIeZ8Jo/QnnYZFBaJdBLmYxd0DDtUzTCvE1luqCGycwsfMWOVPp5bKx281D9GBNBqEwtmhIOz
rMybpUXNh8Tp55R4+qC3OOtdn3af/owKsIcUaaJBskLDKHqQ4GjEp7jh9Sm1tf7soj2ZajE1u7dO
AnzoGeCOuBZGraVT5s2wW6RZD1lJAANftwv5EYTJcGmWuwIkk0f129zhshc58A2L25UoBO4wcz9z
3LvXEkpLBTSfpC/X+FFEoehnh1VO4IclektSy7GEmoFwpUndxhokBQQy+Aw1peUJuFP1i77QCqmr
95rJ8nuD17uMQhH7C1HBSM3oM3x7QTPVgZOhOvRORSCDfA7kb3yl4V8URU0HTxfvg3Kg46LlWuQI
tClfFvJjiv03Ec1g46WNUyusvylmzYVf4wZnSP2Kh4v65ODQlkLWhjQT2G5sAz0N9rvnYoJwrsbv
0/BRF9q5jEdOnlDbd4I2rsjyZzbG9W9CpNi/gtfXSCbEohaAOWVZc2flCZS3uiZLKlh+nooP/uKG
GhWJs8mjXYPzTDaiaOkuDzppWvqi32V6fst269q6taBDV93Etbau2NeufwQf2nqT/ZJbiPxwxGOx
8+7npQ0P3NS36ra9zFU8L7yoPJ9/GdCxCm665M4UMcvTODzL9OkjUX7HqKxBx796zbCwWUHX3tuv
mXByQopneP8rdDGX5tDXxA3miiukHPoTUB8CVRIzRHlzUYZ775PvAXZ5P64bmDD7hSgWB0/bc9/z
dkB2znabd+ZTr7nUMnPe6Dwi2q/zMke0geVJWAngeYdKQBp4mrG9hwbykhGSIArPSBZzqJxD/hJR
f+mrn3kSbrZ2IfFNS0FsFKaH5VrrbfWyKKE4+34COdPACB3CG2sBYrCEFQGvE8EjxUla7SoG/f+8
qlSuYgBpF8MrlZSdT+LoI9NsDX9h6IepbunyoqwSSYt4L/pj75CLC18IWW5znuomohMFT+LWEKw+
5XF7QaAkD/o4a7QUq6Jwc+GDmxmknEbUAMneCDaRSdAK5Y4teECjFxs0oLBxP9lIonHxayXXEHV9
IzvSmuixbAqmefGd8QYPOWSh471otc9tN33K26BzopNAE8Ep2uVLrxlmeNOSQ6/hJd+PoSR0/fzb
RswAf2fdZqZC6rd2kVujJc/VHLEIGnUK4P2dnPY46TYUeWo/W9nh+GOvLRcBSAzMqaye4iE/VohK
+A2TKOyVSw85xTVw9JG6Z7UN28Q8cVr2iE9eXhMxkYJPPKAlKHnGZoOvzAIp6ikH8/7sbInrRWCH
nFptG+j67Nx2Gx6lEEHyoyIwxGGqcmuLs0N+4HRPyt/ZSTacmROSVRT+6wdhTbMnD0dxewRNv4+2
QTCG5Ss9Xa5ABkWYgg8AryITb1pggLAHdqrR3nLmtc0EmZ7keKAIcNCN/eu/fbN6OZHJD3RBOroW
nlixg/L74bKXUhozHMGeJt6HaSXNZCXPSJFBuj6O/ZW7jLvqhWqVewbDH2LAV4IraqPf8pbysM40
Z8+7bFeIJS7QYoUllBnbciqr+U2nG59qvYWIZuBBElxv5apYK6yg9YQr63oZZF43rFYreZ3eatkF
tm50bQiJO7a59klMZt/tHtb8BWF4dYtlrO+/HrfUM7nR8OGjareISWbLHYR2kcamKazl9H94elE9
/od1TwO0xyJTg6YIKBQPuebSj9RZYGYDawZz2mPY+7tU1lemCn0GeGA6JLPrMhreWLY/WFeIzrML
7bntZ+XmB0kwJqKlKSB0LxwIAcu14vVT60SuVu6rQyFg+lOvTSQ9Cvcm0xQhM5PE6JnFY9lhMeue
qlmmosQosp8RmjQg/yRvY4YSnVQX2jR5A1gnBuLkGVWeYVprKTc2nAMzxEdR3TmGuQxkACcKvrro
mU9gVy+MYM9fB+ecwF16YfDmfNA9vEHl64j9Qipo//b0aEavQrR4+rAa/oBj8eH6I8SfY/5EOhS3
j8BCYdQyByGmJ6nW0IdgIceyNfVwbCbKU2ptDCQDlukLZ1O4IzAf3FiphKokxzUsqfMDq/R5RwiU
//j5K5E8sKmKs2dEenVKPkIgoekexY9PLs+TLIi/Pu0g1mMbY1ZWJXTlhUpoGwZpPMMDAGMAy4bW
NgoQMICwSJ3x9/ScTxI1dTDEiiAfefcbVnN3SG6b7HRLVvKJ9FFOAwckoe8FJZ8d3hP+1JcsD7yu
Ayclk3TW4iySKeIhwwkMjZdsy81q5z5twfni2DoqMY6kbOtUeZlby8UON16y1+glsNR88/YSEpl9
rAQpTi/kg8mYvxySHvBsGJSD2qiZkqk4HbtrT3T/ecmEAPvLGNKl3LaBn5ADN7xvNdJQnQE+gNk5
gIXUIGeQqamNCVR3JzhqYQ5+KgxiehslkVZqSsX6BjrB4qTlzKLICPKp0ePrpdk/LcDkg0Axw+aH
Rh8QtsSW7W5w4mXolJYld+Zn9cf6FiFaSvaml45vEd6AiEOmwkyG5noeA8p3V/hcWA25W5yJXs4M
Y7VUAdIupaFvRh5V9G2Ck4gMbBQuUx5qQK1664pnrtmRfR0k0zXUFMwG4G+7zGx1I9OGnFPDYN9M
6CKmirzUZviYGZORcKojpsUcmSmBlh0EGkMwXAcM3VSPJ0WO3e0jT0pq2p7EGGBakJ+qAge+EsOM
mO/1m+lBbD0ar3KdzGrri3BqF99Mtha/9FJ7+0hD0m7A6Z1mXE5ZnRMfnu8gcOGX8VBCwj158Ec1
OGHBrqunvC4SMtGEqD/ZU4O6GTWIG0cPNFXBsg1CsMzpy7pn0rpc6sYAPgSlE/YA2KX5ee3F7p+R
/FB5zgohNUsLmHETvl4e/6ZxDzaBEpvYQ8Dq+DStGDrocs+06ugs6CnRhmfcICRyN7rCOlCFubWK
5nA5CDLE+e91OtAkI5TIk8+3a1L7sYFS/LPpDO6kAOehfzngcdZKeHSOC0g6MlUEXrW3KhKxDt8E
DjC4PXziEIvQLvEoeWQuRmEohjtLXBFcrbg96rrSaNHpa1t/IBwr+YQSw57KiZqUMv8H3tUVP2RB
iGUBN6Hm5wKiLcanDbnQ+GUkYqO9xAC3spr7yKcRvHuvIRU+yGkzdwQOkWyv9RX/Gs3o7fwyU/Jd
zgpzUm5AYRtyybnfbGVkgWFQd9qThIm4W7YMGW0VhOqb7uAf3crCZxGAMiM0CRU/aJeksOs/pqB5
PDW+INtVYlLSni/j2YgPNEyYXPk/P7yyL30NWC8roHhUEP/UpDUY979libtPsYsOMKyivCNzcQOR
3m9wrXbWEvaPx5nyxRpOF0Odlrobv7LvV+fW9Aq1wdX+WitMNLmh0ugYOpKXxETxxVn/KoUAh383
b4bYYJ6JVf5n8gykOY4VOB/sNz3SozAZ+eyPE9imj0f1hkqkB911A+il/FgQLLQuFgLZNlBOWMdm
8cML2RaLmkRgKW6h8gJwlZVgGjM7El2AT2Tl9IIRN75jv1x8PBQuF7pgFo54kGiuZGOZt79BFIMv
mmq+kHHdD+9UkCi2MXHyA66oqaWgVjqyA227uqBM1QjlUBR67xC0a4BUZ6bs5YDGrEwTy/4MVfur
JvdcDRHvWTHuDoscAiamRhrqvnryg527l4gsz5GCU3A7pNVf2MbPmA4ugWbD/C5vKRMVH6ACZ+bz
iIrHW6djO6m+N9QXjK0TOifrjwneVv/iF20cTSx8VnSE7FIzIeMaY5V4pp4nDlKcT0WgSVr4gOCz
4l5G9gkGAzYQBJ8NlOCoonWmm3epXxH6sMhoYPyIQ9+dbZJQGvew909ddrlD4xQgfQS5hzdfbR5V
s4gJPAYoby3aRtRWynD+KEgaOkRvu8B9FRoFtVs6eZ5vtOLUP8Ipz+8ft6IOYP2SZAL0hjvxpqfH
eYBkM+0ip278M6x/FsyR0G5LkdT6iqR8HG+gloHolafot6nEPfbKOGFec954VOqmN21f2QdoElW/
cjw8tYIy31sSt1NvBrvCIecgSyryLSICsiVNUi4y9Ct61WJ84v8SUwdzLW9dj6UN934mViBOWUlT
EuhhinKu30bGeupNGSy2dVl4yukX8tpt50qxjJIXBI80tsUdBdWDbTrHiAWeTyUaMHwdojznQYBH
sIVNn4CTkRU2xIzs4XAJHusnRAn6ohpeVbH43dgqFlD79WXrl87gDGdEARGOkOgeYsvFXoqe0VLu
hnPz+MtnWEMyXTSym66vZSmyYT1PdeuVRPfKN2qSEQca/L+3DJ1n/mpZZvKDDrsU7KecvahfvOLo
faukz4WAlDR+n3744ei12eF13+625SMr3etF7+DXbSrkvsmMZTT4eZZ+EVBUj/av91gq05ULs9B4
W8JvHprege4t9y2Lu+pSUGzsV1XUp8etLDkD1aWG4846ThJRchiPwiJD2223RBCyoHY4LbRemXy9
qFrxuvqWit7mi4JFOdNgbR3wu7G+aMqKudEnJ5WUNyyfFQdIRTlfMdJ+eWCIuG4w8Jpvb7d7ztTj
RskSugDRj0m/OMxlD6xy7YYT1Kb5NRHqOUENNxMP7hWEj4OS8WKiv0LuhvWVVEzmKLDx1TPO9OeE
2k+z5cr5Ia+wF4R8I2QORNw6TAvjSuldJ2oPFKyAeQkcmxBifDtB/erEOV0xJzzE376gRhuoUmGp
O+KePekXCSIP3xwqbtnPD6tPQaO8zuS9x1beUFY6l1hPojiK1qWzHx+iwU9v9CEm2hCgIFXnP/eH
6Gu7m1cMjU5Yu37tDdz8d4VQMoc+vbvcXLDJTIwIKC2gFUfSdlfvoR0rjoa7V1/lRaVwS6ciBZP2
C7MY6Wov1V2eh58mHkzxmLBOTuO/6gtq83MlpdGRGRNsa2RcxMJpeDWhWSsc67f8kiifM7qfeOl9
8+Izg37OV3w8I+BL/FEvq9CQv3oXFZQjnPZp1vYDt6beBcn/glW5SgJtCIQqSsc3jhO8hb1bRJ5M
N5OjVLsA+83V51M7M4JawIvC7N19z+Q/J6HiDRGSGqngZAW/7nmCuI6mWlotDebCGJHONKNQrim3
ESxIGN0FhqlGTIVkmH94NOW/HJLDvumatAeKK7BcD/e+ZBry59NqjMFhWWV3bJ9wQTssnQ5V6Wd/
uXbd959wOsc31vne5hX+6hrUTbdpXFi99pgu+6gJd2Z3+h9oLfvaF5Lyd0Q3Qunhx+YMXgDsIEr7
Uwlp/kyjPnOKOPeDJgB9u2jS/AXyTP0cKYuDVPsfQF8qAYbQLrNzbhxQpafZquD5c79t3BrzJ567
0B2wZWtLrtzuq9Grt5AQrMa+Xx4OHsygTFxV8dxvpOnfbFfueiC3ka0XxYed2FVYAB+JQcltEsyt
QLIKgCL9gKyDAz5tPd/7ii3sMI82twxRrRuaV1QRepawRIzZQpLpwESe0bRhwDC9AsiUF21ln91L
RqR0E9j8C0Ib+X06tbId28oPVwX+zkNwiJ7sZNnUE7eHdMjKCWabpklSy/7rnUf0VJ12pv+zbu3N
2tCTw9lqSPa835C1mleTYKz2/02NScQZRmfYA1JibBifb6yRglqx14FT1mLb3lMNW2I1yVx3PI7m
2Q9hMnIuHN7UqWFIyXc9RjnnPQO9Haa7cvGiiQgOUfhf4GOv3ox49lHmK7hKOb+ZRRmaff0tXkuS
Dcd5NTV4/UFS+J1tGWrhvGprwuzaBP//TsbXMIOC1vSfFR628p/8oE6ZJIK2PJQexq2DKhbtQvMv
FFFVsVUjJeSzKBR6ncIub6c0AK/p1Sb2XMTB30EBhUr7/U5By2zIpc0rHWfxE4rBBrUtk1DTEupG
zQ2HGIpDNLfXbw9ftc9/0dEVhSQFXYbmI3Bvj4OrR5HjMEI0FBR9EdAa2XaPkDZVuE4v9K0S5qkv
Xdv68R9HdY8/t4NCMH3Jg1lF6hptXp6Vl+HzeUe0za9ElR1beSWVcYVLvxsqW1+c8X5Ow7H//tXT
tISsOJYQu3713HTmMRJCel7/ZMsyKXoPPrnJAvMc4KblJOui/Sb8SY7CN9D4cicV82LCMZzhOuTS
K25+6lqBZ0YM+K6U6NJKnQ/0lm4AtFRFR4IZuzBgkeVR5G+AWRyiRCe143fstYFok0esBbzv0UI4
VkO8qKeaySugYMFYokWV78p+hKJFawp9rsY2yYVrzgbDLV11RKL0gCqTcBsyhuzUZx49TCwxfQd8
6sH/bjKRh7aMse9WpVCDXW9MSPEEH8xyFTPNyIbYvpPiWRoiWteiC6eJzhdeo8PCVkZtVDS/wXxk
uTH331xJAXpCaeS7Cgie2aUyJ4JkxAB/vkF0rCXyLU/hQ7oYIl9uGwj7IUmzakthqnB9WlXN5py2
koH+Iwh6VO0lqt+WRNEfSMtGR65TQYVT1U9EBTkg91LmM3HN0KwlRDC4vxC+h7de2X1KDnoFENtZ
IMd3WlccZSOvzTy0PAvL2TNdvpuQiaa+AVDME2KsNFIoZI0dW9vKGjoeArnqA8LrBCbZpnTkIuvJ
aQcHvB4VmLhjxaHfmMJaWbAH5kujrtVppMgyfaWDfLktVrdHNcuqsCX6lUDltH+L8ctYMfxBBJ4V
FAv4ySX3kUyrpECmzMyem0fjfCOTvCQJHiIAaYjZDzZTb2k7/+51NSlhGtpSpb73SlhU12Yr7iFT
sQRUM5jfNwoBIFw72RoxN7nzc+RJyXrReq4RxmhlBLfBNn5xnDZbsBsr9MAB4SO17fpQ893fFERk
pYD/nEndwCXSFC2JrrI9rh9ywIxbQrHj5ElOiulnI/nxqDYxVA7Ehu9QO8ZTosgqlgikEIUaKJE5
9QfaUbQdt74O4kILJ/gyinDucTPStiva3HrWYm2/zg6H7Imw3MY2eyPVWewQdkEGdU9+2YpF5CGO
SX+skVzQAEUkB8jmz3VLrhonzgj5ewhpqi+8lWZEru09IwTD4Nk9iFY+W5rtBkBT1mCazyLIfuvT
MllcUNpLtOf7hEgT1oWoQKV9ydz59loESIX7tPsjA/Up+8xafuSswEQLhBJYN7gQVDJL/UcUdFvn
vEjA5ra9NfQT0Qlllv/KvkkpxTCDiHuJLkctk9a2DFdZHiqsaLBjLvmXcsilYXS9urFhlIFge8k/
dMbJ/l8QfOVmPAv7SMoyX8B3fD9hjKNdSwdI67F+RRaw2qQ2pKWkVlqkWQKjsv+fonn48Bbulhhv
D5jswL3kAof9fmMXDFLk8OHgmvJbzVGWMNTdT8L1/Xpd8XRSV3ZlGuO2VNwgLob8LQQdE0jBKnt8
qHU0Ay2NswcPN18M6LM6XfHpNz3lQctsvQCZY0k33yN+JEKegK5Aa3glQrszxQPfithaH8ASiyHx
/ryNanjLArlfD9AUfYrzRAl+NP4jaZi+XpP91+bzbedv7maDQSg1PkXtQzad4oQ0yfVWd88XdRMe
4tElLN0fkiluk5w6RLe1Xb4E2E5/8aKYaFbGfnKyGIgUu2oiWabUnItTD+5mPVYQMTD6jqMJUluh
ZNLF7BOl/SMOG0V82JZNp6hC1B5cT6BnkBGKDO0bHPp5khNvSwsdJBSfGy3h4haTlUF3Q3n0xLcq
D/wonOiELsXbxYPCTkg0vYFfbMS9HhaCvw5GYGq7ydVKBaDyfFhUumIXmlVfgTdY2/bENbtuJRQi
jIDF8x7B7gM0SdBQKPubKKSeQGUXfoVzYNuM68n1oezhqgTGS73cLOEuzd+gA+787uPx967zOA9j
oZTnXOpUaAOFoeP7tU1MLg+CoO1F7iptERpUyChuAb+5c9glJ7rNId1JhbfyuV2EzzQO0lHkXvBG
5r2MHDOVKTufq9UbW3plvSBU8Gse/ysmXjY4Hxk7eWfDAG8jKhaeuiHjO+WzXKapTd/MwfCJx3Ad
FN16fXCYfsmX0SKKWnCwllWnYwFs5KIx8eDsCHFXuFppySJRF6rUQpeuQfkDZqYIAcMyCKhSfeau
cD74i5CxLoBRWTEWSbgmeBxb5HK7pamPo+TuPXNzOjjeiKQevbA2tLgAcyYN3vqnYxUKn+GC4TE7
sUyh+JHnNoLbtMlbORWq9dGD32UCeGMCZrQtJaco/p8aQQVb9h2wkwFRxbl4TxTOxV60aYqu/Ema
iMg5uLjmAJup3Bg/kWuN6m0hWINKNZpHfEZ1LGIs9AU7OZCuNUlTNaAucKc1bEYHYNrzr5uboJ0A
i3MAO/I4wrC00fxctEbwZAy04hYjSz0dCfp1fLln3Z+wYRqQ+0paBmMSuTlL0WazPjZmvd2UJ0ep
dkKNA8uDRklc9V7gLQcDINPTMJ+dRkobsgvYN2jGCrOHvUAl2CZ39lrG1HiFbrxu6vPDR07FSMRv
Ousf66RW238y7dG6uSpe+1vR+UIOXnEjFpXjlC1OR9NNPmB93qFpsErtm3+GgmirUBfK7+FQf2TN
299xzN3/358Dt1md9ORUHLxfWpzmGOHaaVeObE5HYtIitV/Dl7DSjCLQx8gMCeUWbS8Vgo94k5SF
0q27ibiDLvVHA/ux5kDY/PGRDdXVJ/p5pHLSekxR1mLvKl6/FMwReLNICFQjbG0fPXVd/G73vEIp
5BDSdGy72omwR3/NlpPxshJ+VHBu9+gFv5GgQsbaiKkkoL1J1DTY2FjmEeLyLPF8sIp0Qx8aWzBU
D1H/obXvrLoWr3lO4SLy1UuK0fSdwkNaBAy813BMpMiZ2PfBz/8a+hVUotysbTrJY+ln1doP4hZM
M09VRMs9QLS9GLbjZ3prgiR5ZVKXJXI2KNeVWN6sOVhmVryxpfTakWEL4Kgs59sdJ89NZrLefAnE
iBTp3kcApQdQKqyTbbCD0JogvPagIhkjyexig3lZw43+44MTSPvcFNECWX0furyqfv2SnMj1tzWB
ec3N0Qp4Qrzp3yTRKczWSdKPbjbx5oOAeRks6ucH670Fj5jkxiNUkZlHE2I+mjNou4VBi+v7gOFA
1U5ydmSvZanqRPVtP+371ITO2jk6MPgNnq1gUjMuyas7D/GsK+B4vdjZqSm+3qvAV8xZl1t9teuT
w1urWG3sHZt5A4cQTcgK0diS2aJmEjCW9Leb/YVj6VemSdcfkrgyscMPyCsItmxFViXD+tANI+/t
AY5Imn+U0rSdPOh2XZxrYi5Sb5P8UE3pzX0R7MpKib/hTgs09rbyon6DjUeT4U2UVPyVuJU55gwl
+6+/f2jzKsR3IZ/BOV4yfU8cYkI83+HMvgz9qCPewexpmeLfwwYJ91zz0oghScYoSyRC2u//g+yq
YZvY1yfpsG2KDaohVOGQnKQLa5am7tXiDqx6C6SDn3xAG95fNd/BqMRARClg+3s6VFad0Epb3KfB
8vsBOqdpzwHYHMfqjfue6+Q9pr/i67MoJv0q1qbS3na4/4QcJXVMcgVht4l5M/GGWXwEoxoFVbVD
s86q873tCfb4Ks1Fr6FUPpH0oRwB9b2jJCYCjFk0Q2GGZw0NAd7EFBWVtwTEXUuxEj/0h4D0qI9/
fxg50jVfDLAHyQ3loXNG33hozCoWpyeysinakcTrSbCVPEbSDjrX8T3a5VxJ9MqoRUyDKRVU6aLA
IOqhCMtjuaLf74eUfD99Lk3M+f8N/zTFOoblGfoMeJbBvcE+bed8LRfnnL3IxbemkQKzx7hiAIOp
W+bv0GhAfaN5oNRKZit3Fqaxe56jM3I3Zqm1qed/3s+MVxYSshcd75OXvwF7QwhtWZ/fo5wiIGP+
YMCIwc2qYpa6uCrdgHwiI4ieBm/AWy3nnhasJ28dIBcztuf8rhaHSCa8yy1mfgMyLMgYOXml2SIx
WyK3vunML/twgMkfaRv3iUJlXEqA0ey4LfUV7bbmK3eWAAnViV9BPRHrlZ9XkiNIvrqs/C6MVbGB
WKk/rxwkJqRj5NuGfOeu2PKng9VwOfbUwjf0rwOx5Y/09EfMK+5CJD825ewHz6hF4E+jLQxyUBHQ
Xj7/6t8EWmklrcUwKpchMA2UDXGfxpMPWIhRQsZlD3wYBYQLKLi0DpEkoUO2lvkxqtraCca2x2re
TYLJTyzd52rIj3C7yEnxA0JjQ+hevpqS0uA5uqqXDYU96X2e81n020kUqh3Or8IEbQh8V4fg3+St
EQGJcYPsCi9qtHBR1Hp9gX6Opa8ObmqLx/PN1e5c4/oqHFR1JZbYpqu5A760xDulosveZ5cVeyq0
SezKyCvmHaFJkohhxr7olHw97fdhOkXbdRiF/EMgfc9zgNCf7Lhyn/lHaZdenqF0PnEztrZiGaHM
YUiWZa5AECGQ4bsIuGMlfnrIh035MxOQvDUHMhoUje3A7w97G0sjmFY1yABADHQ0VT4x253sNRHN
OGp1R6Y10pF7L8drLAb1kKvZNxPB83LmnZpLL26ajhAwaEVA2ibgCeQ+EZOSeTQwTfEj7HPyGJH7
hjszqYb6HTG14DM9JAIyaPNmqVY+dzTG5U6BIc3UcYwY9kQGOrtMsXHSlqK8H0T3uo+bMmU0wj+r
6KuY4MDRqJCiYMF5Ghtx5TD097m3yGrUX3QYtwTWX3BMtRQ7WQXm+EE21yKU+4GkN8iBucHC/U8X
KFSHnZO37O3DHyjmNUEi/FtEz5IHNsWNcymeFzZKtiQ7ZtRkNChsDGNrM/U5uIZaNQdRP5iVdghv
Z7cLnVrwtQ8trUkIYwl9j0y5S7k85Yf9foMs4OACBPe1IuMqvBM5q5+qyB8Ta7mwh9eC6XnhckXa
1jWZVrwsHXt1XPvisHELPZYChUmLc2zKtl5gcVhvHm686v4TkfXJQfS1uFChj3jUZt1jibLawum8
i7sxd++hHouKOL+PJR21XUdYky/0ismvzxvup1HBM+vCGnKns2Q/HtFER+g9thh98c24r0QH1Qd8
yoZeejHppQ/I4Lbrwx5Qd1HUfcvbM2XIKCUJRl1x5azUDFkSNJasp+4CPUZFQuQhpoFLXgx7aEMb
uvY7AviH4ar2/KIrDlbBPRaLCZr+A7zxEQzpfZg21oQ/M5S+ZfDjZta7AynBDxR6pgBwmNbfywEB
dDQP+716Y0XiLgh7QNUnxlzwcTgRCqGazqpmuW1+s/+x4KalK81Na7XsWpC3FaQbolt43ztqWcwW
UpKsAqxNcj92blehbYMGOo8wFTv+WBu6eAFuRsehwLc2HS4PE7I9e17IbK7HbvExcRrtIFXw4Cme
EZGvAaoWoLNHL5wimKkKy+7/wDjIqydKSNcr8RbiB2mMqozGzzk1MzdOYnF2J8wvbymXWrNAKoHp
8v8LZmKF+I12TxlwWmrWfTSxvee46YbJKvdfg76ggKz6tYWSABXaKrL92N2fG6/XB4eMywoIh9YE
S1Pn1r1a+5rO1dkY6unQPG7QEcVuPEDFSDRY2vgzi9dNjRqNLw2pi8KO6ziDZhh3FoRWipytpIfm
fCx/qQSBN7PEAB+MUHxVjfSTkNa8FW1wh2LkKTqXQrCoLlJO7ZGmbeXPHpU73aNDyrGfO8XmuwCL
pkQfJjPQamltdMpGKs2ug2KqqKG+SjxPMfgzxh/NNZUYNBjPGPKzmWhrPCfs7Kov0IrxLftfj7pr
4kNMFd8mUkqI1YVqExt+4YqZ3duitg+5JmZwfD4R3VQB0DpjAN8TO/8FuHA1DRLc13a9Y8UlpGGQ
y/5twPpSgFyJo9onPQVmAzFIVqbG4LlRkHv5mkw/LQKWkvHgGCJnaQzzdvdVbMXcytIgSUhsrARR
dOCGU6V41smAsqKtoR3l0stfdTEmndrX97fm3ZnhoY2lwGZAMDP8c4UIw7Koz1Ke4ZV0cG+IJEVC
07RMfPS8QR6+oqnHryI7AafBs0Xf1xfaVumWNTlqbMG0W/l5YsaLPUkxJAtBrUUAcM21bEwei3Fj
JE5RuzBl4DqJpg1fLuXX8Q7yIcdBmYQ+MnuwIZy5HWJbVhPWKwKbTyQZQJMrubQrk5BS6MSjZDp5
autEm02sB0XMji750d19+hEIsJidZ5Dgd4WD5j2btLXPZrKLAldvPiBjSyqjujIY+hgLy6R+cKj0
EnO+8pnFPwzhRryNty138Ef/tFMyxr6MHUopKQMM097xzHYHGzfU29CFP2UsLP1eAbS05DXSSMZt
hBBjq7D9lmX4GxZdoIWJcmetN4N9JsQOCKT+UrGD5BmHG5FMIZ9KqGlgd61cqR60yDFIf5oWPQm4
2OquS8tLoMhfDbXKEJsz/BhRtEhZ5OUhCkVyXx+Oy/h1heuMJHXhEjeoGkfUwVeaKnzq97MyMDcG
GPVTDHw+aNvJzZDFVxQf/9Wm41AyMeQfgkpNLjL7nuZ7QEDciKEE83weYaAYCm0AAdzm81GKsN8Y
WfQ6p1owmAkCsf47GswmM2CpRbwCQ09QmCRhsNKG62vtk+7ME3yA7VqdMDfOCKf5t7IKsu7BBDVX
gZ33QPLcipcZhfhde7riCVGWQOJh+52ouOIdpPV+HytfHDhdRg1ddb306ouRaAK85fYVlGGkOzwM
eUTRe1SONXUWqAupcs+vNrZnCJTxwjc7cAUlixsKbfXg679TjR4Qn31wwXv3rkaO1YVriCZM+MK/
xscxam0225GEzFhx9JHX8HBL6fpNp4L4cwiUu79UQxqxqYeLV1jK3sze6+qLmAQFHNjeYAuO8YKu
NHpBdx8vflOs7JC5QAcgNhvePO1x//2FI3heJ0mnFCbU3zv7G750yvjI3URCc2IvAxu3aDXRYgX3
Firj3K5GEmY8vVsU6v77lz3BoR0hRMclvlEoN0Zx5JsVb7yLo8QmrhYLszjrHObrnRo4cvsqQgVM
GCL3p5dpXSVLg3zPNSuAfkwsqCIjPxKwagtIq43a1X3Gv4PyMZORCCyqCgdx+DSnGMcHkhudJyj4
yXpAvoOhkQOvN8LfkUyFNDWStcGpPKf4Kw5Bd7Lcn8mQYSUZskhSwC6va6VcYYTW7Jq9eDAAq64e
fMHUmoJYJ8mGEJq60Db9eIeRMDOLNVRbb3IVLqCBXrO2LGt14sKYwl/e/5qGqJOgAyIflHDCam5z
2BSS2yOxzT4yzpzNi+T5k64aUL0jRYNYV5rC/ne6X6LLY/txEsLSrKXDhcmIMHHk9GlDtD3Cs2R3
/M0HAvgPK2EwiUIOyrkCd/uU4jcqHLanrBtzSXtresxBP3gRRF8/7LvU87/9Kha4nQzraeh+ebq7
vSngQkHCBARJ+n0VPjzFHHTqPQvLeCYQqcYacWih6Ka+Xk/beU6khAjnAUECO5sfcne7WH2fUqPq
MFfnO3M8RYx05KvsIFi5mZOl3YBfq+9myn9g2y+yJGGnqfLydTywpCN+PSMjryOUZUvGFq61vv9l
UUUTcPMjVdYmZzMuP6Pp8vokM7Sj3mUWE8NiGbPZ+3bEC/SlKHRe4EwXZK18MfRrxAjXRGxFoIri
Aqk+Bq8I9SpJWslmNHs7pESbwMsGfsWAVKdJxU8f0wO9NOYBsi5kumCaaVEduLxzhBEpIB6xI99R
jYtCA6uKOFvzILPpOsl0z6tL/cIc0P1sgQGaDHHtq0d3Wz8UETG1hYrH47+UChIzH4IPPMpxa984
VO2bXMMpFD7gf5CDqfWp86QtOaUyRVap7NRPKbV6IGfjCTfyLxWccwrnE30bQ+Ka4/F2oYQ//moD
CddL2035uJnoDibW8f97KKcTkezjHgCtbrGKc48wlZkfWCKeQL5FyGpLMPnwTmdRan5v/OFLPuxo
NGUtEfUdg36Ncv38quHl+URf5WwPguoIgYA87fmptj5d3Ifbi4YkkKLU3awfGs95xm/1nF4X2tzX
Y9ObjQWQLh5h6P7pUG6f5VXXZf67joyynO3pSOXBgIhIMidmlr59/NPcgARxM/FJf9i2zkCoAQ6z
jtuu0BSCt5wgQVg2lHb3/Y4862PiRZfSBytG9yp4RW0AiKIgH8OGH0lCDJ0Tu82wl2m66AzqHp6t
rLDX2tA1cT+jK38Dx0UnQV19dUbYsOAv9f6FPTH2Wko2xTkt8m4CcWyZcjly7ZXn4Zz032CrYMtN
FCh9j4H78Gs2gAntVnVRnowvJEuGuzYRtMzhOJ+bTlkdb0i4qUx2N+FiXELoacc3dL6RvkSc11OB
WCRuvjdkeYEjotpgRztHx4knzxazRrhbwQm6N8qLVSG8q78SnaqJL/rQqW6ZsO+/Pj6WCZtaamJp
cBFc5d3nK4qtVbzWO0u0TrUsHRU+/0nT11MdbjgpJBvkSLzWu/H3WlZoK0ysh5cLzvIdSYrk3Pg+
CSeQO2C6xxv46cyna91g0ZgIcTo85qV1gulKV+076Ynk1FC9eVNeWAeXWAJkLJYk1O3mhraTa7ae
5J8bGGZ7bmCvc3el5ZeKS2aKYl58WtvNuHCt5MeizMt6GtNP5eHkccQ61uRkd26KvvVr2nHixhbU
w6iRmy6ZJ9v0rZ7kM2S7Eckvju2ncv0sQocWll2c3Xc5eIE649xnJCGiQxPqWeHEcLNfKi0niorQ
zzkK0QZL3VLSeKKjcakEjCJ9S6DDDN8QL+5H5fLGa2+WqGbmF5irDxZKB1LEWaoSbAnPQrJ1nYcj
690KXRZNWEeYCNZDusljWcjV26+GXUHDDguXzC3RPhoat3WaRMg5VGHe8Ron/tCeQhEVkdcZ0ZoO
j5Xc2MvU9dc98dVCYIHf2M9kL2arIBlmVw2I9qawqpiyttUHsa+luRPeVDzGEUZIkLctC6QkKT7G
XexDCTL/8Yvo+urW69lDCB5istgCluOqBpRA520Ced9lbaPQnC+KK9OqfJhZOtipOlTOnIJnG7vp
b4JeQWQVyofXFEqN8fWZgxpZvLy9G8yw2Jtpnj0S7AHrL8WWfQ9lEpT2V2DNW0uynSoANZknnEh9
XxjRAGWV1U26/xHkAi1tMr+HFXcttK94wVo7G19NNMBa8c8QTRkiHL4k0A3pWicuvAU+q6ygFXRu
2oWUeLh2rWXlR3q2ybfUvQbrWWqrnVF0R6eN3ZQ4sTFwjFFUqUOjelV660GbcBD2Lz1JGPWLXEt2
v5PNGwMYwdqIuVITv/eqW/qSHqD4UwhFwMN/7pzOxPZS6kxj7Hcho5Lo69EqqJgfiLc8NhmugOS6
aAxssUSz+8ibkNcTKbdIB/5w/ECQcJuxReAECOtEJwlNo1oL1183uO7RbQJYNE4MNXRDZ8/CYl1t
DcTyTaWpsaO97k4JJTJ/I71hsNktRPs2n+Z/X8Xf/TvcBJSMrmtGRWJ4poi5FBNNiBdurKZREulJ
W1V0sX3TA97XfxPVUpF2A6IFHpbRH1cY2486Gjhg+4yyZ6v1enl9Eh6dpdQewWXFOKMBULtkYPBV
DbTvDw+lG/uN43QID9zOEjPTKg6HQCy7TDhjJOmWDyl5aSs7lfThVASP7BmTeldwcIA/PqKgzTm2
4ACJB5TY2Ajlbj0QbG3bmhzeQ6hp/peHxjuboTsYYKEJr8RcwDnq6vlRQIjuzEC4R2hvcWsy8ekM
ipAMcCaL7Tx5eODq3lvM5RNi3QxKZUT7gfSGgyVplvnPdek3SCfioMBhNN+lVbB26ES+Ocik2sgo
Ovn4hXbe6TE0WWQrSFIsO7hJioJI4JGvybKmeoyVSe/SBr4z4QGF8d1IZ0mOTgUysfaC8RwjAsxe
qFV3Dr0jBwradcBb7vPiGoYsvCpLyBjVNgSGQJT0Uq30/lxMcWXEpF5X2rgdBqAgsD64tk3HvkFX
YFnK1fjpjMDu10UMfduqebuk+LZfooZGrDXX87cXtJXVR5k0RZZWHs2jQ7b2PEVa4It5wR21XXhQ
Umo7ssfrniyO3mhEMjke9h8O2QDmar+kx5Uf0Y+cpI9b1aoNOhMWnqZK1qaqijxhptW2drIjw6N5
t7MeRSvNqbl8isKZPmJm5/A7/oyilqHhy54ZwYVLPEwlaoFi/jFK26BE3EW35dmVDnvFuHWrSuCQ
VgDtz4aCDcWB3Ysjqbm03Zm4qXcYr2UAg2KN3YFSwO7VOC9chC425BB54025dgyhbvb0MxhBXC5B
mg2Usokp8XaUMdkhch42wmOiE+UF2Pq2HVKN0SAjl5RHl3Z/AwqdxGuf8aVUuGZgeTp7RpQ62sx3
MZqg2q6+DDKyjt2Og496x60dYOUoKUQ4z/G6nNEmiN4pP8bIh22GgdHG3WCHzBSejFhMxtoyjNyn
j3RAYOfArKxcHb50DZF0FYNA2mej+YXbbwIGuQ8h1mqelr+XjGXo2LVY2Fg64QLixzU0dBO/5vU+
PuXcraoqtFxwbZldjk10hBhy5+eJub+f8RvCOazjWL0gvYpsZns+3Z1qg/79DGQp2T8ANxcoeD+K
jdpZeJZrcVxhhkuLEBmAAqV0SrsWaASlrWEilVK+T2dZ8yG+bM7RmCZMVSDGQ+fVdd236AQtKvBg
Vr2eEAmD8SmECvNVoXIMmM9yZzzY4FZRIloNee2kaifsLcKt5YwikRDaYYo2HokqtLXBdiDFG4LV
c2e5LjOy97qLSAGDDMdKd4KxyiCo2+X//p4WpuehUD5IHT5cy2iUIVOkuWljHB1uklkVw8gv7NKu
tULj3lEJQg8aaXZCO3AMyulv6zt8f7QIvLG4e5NoFwlOKvgtAs2euIf+jTcvEuo2HH6V4TLDrgMK
36R75eZdNNFn0GOYLs7+BAyt6tiexrswIhRBLWOGvF3UIU0dsHxzAgiQWaV3+3cefyVqZ+eNs/dS
5LlDgHytCvkb4EF6O4aIyTjX3293gVsHt9r7qjdBoNied9/LbnjDXh7IDgywwgc6hvL1nkrLlKT/
7lEs4TLta9zqgvb4BMCUF6z07wlTTm6sns4Ari7u4Rlo/6BYp+mi1BJHZ7ZrhM3hr3mH3mKlmSEp
gsQ5HhkBm08EPioUaGWK9LOcA4l0NsjdydGB2Le7fJun3i6p0E7VVtZi1WkrTEFVGe5UnDgL+Bu5
s3ZaVieiC0QI3BEIYxuWvPoNOhGyzS1BCinIEV9jW44g3nAvNqKDzrk6yVRX5xC9gHU4Eqi13NKV
QG0RJxapaYUTz+DBmcst8KOnuoZnChzd0YElPdCP4c2DvtHOSApEZwWTP05Wz5mYkvIXOibUzm1B
tOtpMw7k1pcVM3IhaIskp8FEyza3HyvnOxkdeSPaZuWSpaMssE9X5AvncmKWCb7lX5c+zfRTP4Zu
EsqbvSF9LQ6J+dc4FKp16aQo2aW78Hzzxpf48EAmP2afPr4niDOO5ued+OVbW7yCp7axjAV3M5Ne
b6B/TOFWfpnwSN4bRIcXwS/jZxsL1H7PlCXOseSMQ+qVf47HRRUhdWEyMG1WzqEZPkqDBlOrCdeo
66ckqxHpcxQsGqFLRjqvIMvAG6wnpjnjFguoU+kSS6slLVBY3wOgkqEYXyhhRpN1WhZ/xXGvnWkV
i8Jcc9a2VYQJJ2xWLGmCRnEtL8mSPaSgYab5/HyT1/skaZJY5KLKkHUD2qVYTZgpoGud751fZ284
GDrjoSDj8yvQW89faGC+dhgg20PfZm5FplEiikezPfw5PNBHZM1yQKM3KSVzZJlerbnDSPXX6WZU
2xcSqHPdTzRllbMxhNLa6rVdMyGVlRu5Pxe3S4cfrKNfYZdlQiAoMkt3J1oOIX4a0gU5pHjrqcR8
CGvvd5QnznvW06vpUNlIOTwGBTsa5aPYFoy1/KsqRsujftUspO1UiOIwo/+3qUKcf6gfjhQST24d
DmZYCCYmSR16PL5IGZF7omp+0iiWVLX7bfMwxsDEfKQoZAK55N4IYJIiy0IvNehbZo0Nj74o3ylO
e0IN4ai4/lDUkzWNnm+kqKWYm2WuzJgLt6oTyFpFDAQvBxs768o9UdPGPvlGkicC9NFbnOQcdDTA
KUYJQwqGFoxjT8NJ6z844r9SrnC0DT6admcisH9N6VquFydnlJARdwsL3nKDsiuqYSy17XIKOC30
R7gzrpjWRe4cenXOeR0wFczFuumFhh3zA9sFQs65qov7o7sO8pYRq2IfvVqH6wmaKNMf6dKIJrCm
/hWvKrgGiQXOQL5ifTmiCZpSF7yn8pqPEr/MUXR0sZ/l8kyuJVkEWuojEP+yFDH3X3QSduCmtmGL
SbmuwsKwJeL/BmSh8Gs5KKp3CbE7dRZ8fbEz/LZHb3c6iGx7ANs2owmEzlGcqDizTho6/TMVorFJ
asjUGbOw9IeL12GxnoldFg62m17p2CpU5dJt5LlRMGX/IWcdzkSRDYqtOxf5Sdrx0TyC6o7icQ2l
wS0BGgoKCdNIrJcoRCJWmaWhfHO66b3A+/qi+8Kou2PAAU5zCKT5O8KxMU+8bii36OpNB1ynqxnK
83ZfcvPJYDraFXdonXIckqAnmMJEKzNbtYeXEGVsP1dNtfA5Io2sgJzxuE7+7gyPusX2UKuhy6n4
jGhUIeyxty5EhXwf0qccvI4QFrF3VAObUpL2W/gGzRiwkeBohPFFXN5H5C1EpHC2/cs1Kv6oTwFq
kCYRMO3PFbq67fSWH5USCWot6YcXdhsObDk4zEMKeWYI59AbEOdW3peFl73ogHM1bsF488HVTpr5
SgeO/aGLn55X879B6LaDZTwHnASQ1Pklcm+IztVuYzSw0FiQzJE2lvjf9XTiJAtxBnKFiAu8KbFu
B8CZd9+3i37kTt8MJVvlxUI/ru3XHFtmO5yy+Jn79FzArJmPq59MXTt3MnPReGrMuZ9DcLJTBPFH
kf0pdQFP+047Oh+wTsfJmuMij7fLDTknQ1OsJl41EO39LdgKCHd3hKndS6aAozAQEvxphQ5UUo14
YYOK5uxc1eAZmT6eUtdR9OSVVeShpzMqkQYUHBCqMk6bZgPAAltcDhy1IXM9p7h/CxAl/rr6JdMe
bz2QQXLiIcLQTeXpj6JUo5OAnNVb/utn2Fsm964DpulLP3401qoxTG2Mwh2gaL5uenErizomCAVN
dw43GYrckuqcV2LJlxY+JMYbhn+8c5Ln17QKbY+38IRujcEgtwhCj1Rqenj7WAwY9IIDPWZHgWWD
EnRVUoSlcQpHnxs6pY8ONrwBl/yvAgknrIdUe6dsbpnEw/GM7ZR3Zy61Rn587O6jFhcNxCF/SeGf
xkwDJWBJJHcAXW88AAZ5HSSUzwM6Is0k3ldibq5zHuhQi4q7rxX9j33nbrFCYt1AjJOaSSgj0spg
3WR2s8ERAsqrvjq9//iDtSyQIXwzlK+gxKD9MwfRDWY5k891hsRRaxb0EmzuON2qsirREkBCDxZU
WfJ50cgSFftx9q0D0gyCUEvT1WGsynCDZdPOFbRjr2u9Zi8eUK72PENDC9mi2NizVrt/zJteWo6y
UZpouEixsHvNkBO4Y3WyUKgm+povq7qOX76o8HkVs7wA2x4OyMShNbKkvj3DS2CCZtfSPWFV9VAA
mz5ZAV0m49Es9iNPZy4yAFvckiarMyqA0MCnJqp6Aoj8jfUhqbi+iuuguoWlWGQImbNQKSKzEbOG
XRwjl8MQ8ov9kF++C6cfsdg4rgQCX14DUD7jQgOzF+cvkgpXoNBInNVoy8u+1u9JsinZoEZzKhNH
b0Y+1gQgZpeFjONGM6UIXI6HO4qHysJUP7FQ+pFOb09E+ldzbEeRriE2tCH29LZqQoSGRGe+suP2
oktq5u0WL2oPwjf9JuEWOBswZPcE7eyGwmY1NniA8Wyh/yuuvnjkHUZxQRuJd9Im/xcNf3pX6tC9
piUAvKFcmBf2417VYiNSZ1OygQG/2Y+u8uDfTBo5eENv5w7OSpRNKFEybaoeH2FvaeaiEeXBPfA3
81q3lJhCo9yTTttboMz1FmTGqiRxe3m0QQjIAC0C/u45cb/TldQ87zYs/YRAmgqxVieUWNhv/pTZ
aNJXaPcAV0jTGKAkpePlXbs3i/Bklt95UxEpmAVvEhJiodHzinDOmeqJtCnDrdu1ATgIHqJblLx1
DGPRvYDsVC7/HYZlcqH5e26PVAE3JA/2W/tN+BvLAWQXyN+llRwyKwyAQkrQEY4wfdHlqCkC2Ktd
tMaIpIrfzjE+6rvmHkC7r4GMzJXV53C8U+tZzU4j+pfSiLGGs+8RfznL4z/nky7ovJ+x99RZSW/x
UHY07daKDiB6NLv2GFCfnHloXLSDy5bQLVP1/FWgdV4GAmuE8u/aApsm/2C/xAQX7xFYZcAP/sTk
18gDzfoA3Jdj+AXOJqx7x9HW4xSCaFWI0kmvMGSR0Nuhz8bVfQ9nacwgRcLS/dhEFuKy44BMD1S7
K04DpCc/v0xjVqeTEwDZAj8GwdQJRfAG3jLnVsvy5K/Y1M1X4OaKeoY2VvBXAOFDso1Tdj+E6Esy
AZxOm4p69cZZrjdGu2gGp7AcbWQ6uRVciFeoHBKobANFEUy9fLG1ZaWsfsHhkxMvHhOHo0SQzbpt
dnZbqrydwG2xjGFBAvwAgcJiQdv40yxxGGhSubs9kK7pkl7Efh1657D+yJSBGOdgy2ioWEZVMfUz
IqwnnMuGvkAmAmOduQG3V1Q5wzuuYWyEYFL7GoKYxhxsLdhBCiPctXVe3Dbb5ZwebgjD4kSpfO9e
JjKW/V19VDR82Y6D+N3qDSpZc7EmgXPR251+Kvp/zEjebwg+WQNgW1HQ4MAr3rXZsB7NnsyZ/W3H
zRaXihKs7E78Li+GqJ5dF2NeyMZeVfKEkp4dAW6EoYmLjIZhhuoP1ygSS9tmH9OXdoeymqahOuNx
L+kf+7EGFt7HLnUOkdejRH4RqvLGT8vfrO/cEofa0rrOM3lv3KQVcvYSaycjCVUOSRgqqSeylcaH
1lIskH88MSJeMFNQOuCzTY0EpvUzUTiK25Hs3J4XF8xbJO4iFCYNZmgUmYXbxkOsnEdptliRkERq
EN+awN2iEfCo7/esDR7ahRNmpKgtKb2dacelLgeQTphND2C0Qrat5pBwL2731pV3oyK0yA5uGHGe
M99AvfaRgXYdMymW6o4VD0lJkskY1Bp6GUkWYsbWHP8Xxm3+Vp5tIkgzrW/iuwKZWvf7tt1+xsGl
tidD7kxVJ7+3k75wNvMJ6qWMiqLVx0q7/Qc4tt1G2vu6V8hfo8xrm3wQsxKkiQhKNhnHn1hUwZ5B
qf1NBpIIDsKRIvTtV2gxR9RfLlrUH30dFt7LUrmUQ3Ok5wCTiCMFysnyipaqb2VeNAnVO7vvzVuR
U5nvxPZaswx65jseDuV9B1VTxTFQ8uyfPQKudeZQqJQyBZHl0K/wD5s2rFfmc+qGMDfBzM6V6YlO
eBe500YFrVOBY5S0c3HeH/xgzWVSp50e4/ZqAkCl42kuVEJXY1vdmBZEkl8H8tVmy1NwHgkkefYl
JUzQTdVjNxZi5YfRbba4/qGo0XOa/3X6p/UB8eg69+irBzmkD53XPYsY+RFXFRSP7FOeGP1M0Fxb
h5NoD3M65EOM8WjUAeSWYS31nhlsrXVqrWVr9viB88GuFcfxeB79zQZzChyECLZBFfqDXJQnKRCk
ApQR9eUuQAt7tzdsmzwjrgtlhWlF5oMrfDtxvDRt9SI2GzymUhLdS6AMq7RsWM11j7HGi+Cb8br2
ZlpGaAzXoEpS9bpiguk93ZKNJ3L8+K+hH3cDXUHS4ar3Kj88hSvVTgDRI109Dik1RTC4fb2QEdQR
QhRrznTc8cmwJjVKZIb93rMXwILStDJIMgIYzh+d+6RLOz1f3+GRBqsqFKgoK6ae1aiv39nU1LY1
NpCxE1pBiVgyF+rj8QR0ul65ce5Zp8Prztyi0964AEZBLG6i/N6vGjBZtq5z0pd3SGlbav+Fh501
slEGhtimz/6vMJnkP0zJ14MsW16oEg2HBYUg0L6I/BK/zLsCGyOM7RjgN2n+uo2hvCl4++LVZV0q
dSEmEKoU7QacNcskZM5SS8PzPmCkTfQDrecoe0tYs+RR3z0vUCwWSepMtcrC7lmhNfqxsQZzTWKy
l3iQy4DjuwQ+e5r6FRmihHM8eKywAs/LmyoglYlRedFSkGsfdr7OapqwA5b1dLDqaOIKE41tsXoT
MkA16CTNyf0JWaxIjQAioKnv03/4U2PpRRxSHBjcLx1MV14UMWP5Exah5qMxd3AUuwUgAhYUwXB1
WtzV0+e0Y1u7RbCGvjXA3aqg2Ag0FcIaeOm53noIoXHp/C2VtONOgjrxPASodWj8OJ7jf8nkgswz
We7QlA1yM90D90Dm9XAbRArHbLkF9oIXCZ+G6G4fah0TW+omCq4MKVgPUYa/40FUt7r4mwNcV9ob
xrwwgR/4hUcyYFKyR/x3Kx1Gq2YpqWaFlUR9138CknmaG8Qupwqr5YDbYFRxNG2a5mqWmwdv/VhP
APa0W442fIM8QDN4sY53Y35bEVIjAWLGcIvlQ7LsZAQOOTvfFtbM6GRB88c4femVFO2lyCaR8XlJ
2CyZJn3LIzZGWBPgP7to+v3+dh9KDHwzPlGoJ8LYlqQg2vc1Gqr8lQFlvQ9th0c2kYdaBXtCkAlz
gmieb+prj1oyGNGhUnamgKXF0PIWQ35Jdu1fSSjJlAeYfecOtRuvtE/zfJo5pUZBgo9mABtW9eXT
ur0/il2l2x5JDlJ9454AGk1SfglRtg5XyZjlM7jDDtY+sXTdoCThJvUBBkarERRQp8q3jcqLTcUX
ff9EzZ2ggeiAW0pUPq2lBks0MSen9o9CvVFYPnvM0Hw1ERdPubiIamFrXJeyOiUhUEhwGUXj9U6h
wvWyxMEpCJjfwOzpsz00gWNwroA6ZUeZxfTn6WwCRI/RJ2p/uz3oUJ79A2KHh7uxRp4hGL+yZUsX
tL8M53AMRtfFcSUXLLJ1gBIkpdc+QeXUytb81zQcd/m6vxRh9r0srBGkkLPBJwbonE65KSIplOkJ
ZK0rRgjv9wn5XvS5Rm2moe2q9KwJyWzABew1gfKvusPv71vXDqjQTHYkD0U5nG/vIhuOpjohuCCn
w0NYZ5IvpkXKRQDmc1WCjQyy1T+Ruo29sI5kC9MT2hInLrV9Xv1mi+dFE4T6CqNuGToFrEcMqM+i
7ZVtiBgueznc1nyZwgfszya4rsu5J1MMC2n/pU75IJNAuggsWYp9YH8US9OpedAkiXvmsyMlN1oR
ZD7m0gmwM0qrNlGdZJ2fVbY8OdHYwG9AoB/1B/+936Xj/XcFDes013vfbTBrHUnxKa0hlFrp6r+G
5g9M3whtcOuw67DuKyKdeeL/W6PJ3m1UPyYm6z3qvjuRvE6DdhGPkQ1DRz7+/CKiK57IPucJRWNx
D+ezYvV4yMoEDcU12WbvudHekYxyrMOBcWApkqij54mXbBmjU2CEgfRa0Rm0QRucUbU6L05uXkVK
lRGYPkqfhmxEh2cl9b493+zs8ZICX3twLoiYjcqtICaByIrI+jd/GH2WhT2FKSS7rtiPSTtD1U8V
gVsRBgFiUhv1p1wvkorAssy2L6hDQmVFgeRS7MPm1WF6FixNDI4T4Fa6fo5MrUkwGgX9eazscoaW
o7jnN+3DpTREnBM7nfk+2d/CKZidvMSB6A74UyxFkPKGjuPnM47p5Tm7ymkUgzAfnyEDaX0Qf7qO
wysqDa8GPcBuofM4bM07JS/dRjC8Nk72biv9k43IU8qb/TRppGXKc3j3JesaqeI4ZrjAfqP7WT5G
uMd42LDcpI7xYtsCeZkmSLh01+/sK45zhXutBx80pk8iRMSQXGvr835XilwXzWL98seBBK8u3LxV
UQ/vB1QjhzYwJ7Hxsgff47j9zjMUxVOAVEFbfCv0TCtLQVidfOeAS5UwQTYOLL/CevEBVF0DeEvu
07GsSRa8a2KwsSBy8u7VJlkWRjknQKYJfU8ANOCCpR7BlZe7oINkamh2/kD8e0xeaqm2Gvunn30L
5qq8A5A3RDD8t+dAeMukS3YLeOrQSZ/crUlrsgMlkHvvCTBu8C3FC2gLe+KI5w3AtCJ/NMpjQKFc
sxuNvi46xnl6Azxn2hW4ewCgb2rgLwqWDx4PO0ccfqoADw1pzb9PVd1MxkcYvMaVNrUda57rKggD
1WKe57Gv8PI7RNg/kKVQZ8bRxYQH+qPF/9q1emKj4BN9jQxCb472++AhvTCEyqmJsSAyis3+3HQ3
7WbfNqrwbU2vYzlm1iuRUthRCleqbRzNQX2w7t+EAI1ZgstxE45Qm8Zm6L12+eNtBK7BWdOFgAe3
fphEPIBOLt0Wop2oZtGf8GzfA24ROx1VMacrIelZYMyUPDWHh9KrNzrejRQTA/pCt8E6COAJ3EFC
3EbOCLIF+CUHXe6u5kgUe1T2EIDsk/vqGISv0t2H1Dy96BGwTon9xbIXPPTYRUgGMlCAVWVUwxMA
LFPy0Be4pAjLmpXUCTv/O7wgY1TygwjRehBubfRlr+NJpjGnc9sIhGWkCHPtswRtRFOwQ74L3egs
ju3P9d5v0ut6v9eAJuv2C4cOvzJA+s2Q2slfDMrUaZwxnd1a/+g9zWqGSxMFuLj1IftKtdExd3PK
VknNJZyCsr2ZVTEo86Tb0fA1lgkObRPiqiWrRbh5siiW6SHkOJqjtN8k2qdROPhNvuO9ICmYmAES
fRiYV3RLIL8sEJ5GXpOxH7734zt8Be60TLkOOmnWQZQeEuQEzRa90euJxB0UBFBwbfMSOu8OV4lj
z2M7pQaWTUJ41nGt0N/5mdxQbg3hmcdtJ2t0+dgXVoEJjdWB1Se8hgD0pX5hcpNCxhMGV9jW2o4f
uGB7ZNgaxHQ3cojTPre1Y02HYbOngR01Mt22PdMQbcHtkeLT0Wv8YPNGVbrS2RRrwRM6E2YdWpNq
4I8ZrmgwTZqe1a3xXAu5M17QnRJZPCYEU/JpQEAquj7u3q6a0UVIspHm+lBPnMXZG6J+NUfcGvrs
WTtobZt3mbKdsIqKMCwtY8d+TAC6d/LTiWe5RQZYWHqclxB6I5n/Gf+wJK8ZBn8JhqVAXrx3THJj
WznV3jaCaD2abrBJxjALA5lZXW9Hu8RMxRFm0HCZwtNQzUtOUDB9z4vTnwLm3dzhdQmv0GbyyXdQ
geWSt5+ad9aJqIWV9faPcvf05fvOMv08SeeE4HrDNC6ft04+boEX6vH0Csol4JuVdbd3tfVhknfB
lV8G3bLotOU4HhBZHVzUOXQbuNIquHKM+1nXm2nSJ3zI8nyGyRIYH7x8qII0q2bqe203vU7VxPlJ
ZfkWR0X0f0TVnqwLc47uKOsJxN9bWFigABe+o9YEWwouA0RUYixmL/cF5PduwyUnovKdXB+TvK/l
w4OjDdfKn40BnzCXIvO4np8GpkU07KSRmmCxP2xkD5RBTPTFard4Kh64jpbPELeEBD0vC/KcqVEG
aePOKBA4BCGHTKugu2NZns+NQ37ibx/OX+sn1+sltHrGr8BqC0Z5/rexBAP1HMGMTK0+pol919Lx
RrNTM664Vu+kSLW03fzLFiPGmOZZC52044NMJCCovVOQIGBC4673xar34vnz2UbkunYx8vXkl6K8
LzdlNUYN8fM7DKizpn9nEt9/rhYeklmZ4d5ilWdaMEsUOQ65/6uyhffGuzSUbvpzXVpNdxWtaEXY
QFtndK3MT+j3k7lBu5W9c+CsSao17uZqWm8aMeykbGJGdktZcj8nLUSrYHgvtLCQFAvbmJvDHFIT
LZerBf9HQsK9aowojjNPldoVVsGG3DdL9uNVUDdXv6ZMxEYabeEwRgFvf/WW56w465FdJNgV+/b7
+Yyz5XzwjWbHhHxNHLsOQGKSIY0wsJmYux56jRJMyjw0R0F6eNpUmDiuUZXPoxq89YPhR7mGuFxA
fe3gDttVfSNNaIS13mJziCyr/sos/m4BxRb5pO1nA9wh/S/3Phc4CE7/ZZRH+ljxn6SF+B+YYuB2
MbXysaEVAFOzXOSUyCiPSQv58Qmz/5UgkhUg+T77TKz8nsyYSLcXqyKGA16dGD2dRCQCBWwLwXtN
Avrf/3ODl+Bz6oeJusMhoyS/2HU9tDKFZQN1GI8tlASnLhnUykRYtZxywtUSHfzol57ErStJdhJu
I2vt+3UOgfGQU99Le8sUK8UbD1R1jRMAYFAFADZLQ9op+qhVg4dpE7NMNrBu4B0qIVNrvyDT9uGj
mOfRc+i7TIaNZcqkK+n9aM2HIS4hLzBkTFKugPokLcD3yIGbzU7N4UP/HOoBC/2VLO1Wftl9rN7h
Wsm81oKXVKn12UPrTqXNXRi4hwB0QhXDEnzuDW3cGQjbTPg0FN2zHeRwmoEOPTHdduIfU9ZcxAy2
cTIxQkNCrp55QS+inNh6RZnHVRRY6ZXuAv5aK5H0/RKx1EcUzfILSBsMTjnPLgkIEqcxsJSAOx3t
LIUhLhb/FtiR+3QRvcHVoUXuiOk+YjuqVWbek8WWP84hl/OSPBmeva8ZrCMkoyfAg1atRuaf3kcB
P7/8zPeuYvXOYJwJhbntSw//BO/ydM9W3lEMzo1bUqt2+A4V+8XqnVASTmJJsmt73B9en9UZ8zkA
pIlsuS+XEiG12MYYZTIbcA+1K8pQ1t7g96hgVto6DoMoAbtitpUBldOb3A3sIDzdSwTrIFR7vcUo
vwohRW2cZAZbDeF6WHnL+QqeRc+hUFW8DLsDKLc1ZAi7S5mUAxcmolqRoeJAL46HU9qBYQ+xUlcK
X2bXu/Op0pdIaaPYX9dYduHSlLjz6PyGQcAKlnnWeTiNGa1ru5w1EBqprMhgGWnM0DNeSLSEIUBL
pE5OfIlXE3LN59E433tQk0Uei2a5F8a4Uikw9CCnNSziP1l6Ijz0GffZmR6J2X1rPZfaYHcd8jBP
ZoFbae5sv5YN1yKp5/mwZQWof0k4NUnHSsrYUIkWCuxRU3oMG7KRBdRNaJPnu1fKF64ayeiu3LeA
C/3/i2pXiylDoTawXTPkZKXpgjZCgYxAob2eELLrrmMm47fx97lGnAoPJf9CwrjwBuSKKqe/m/bk
wUfmxpGuzTO/Pcq3fF+5oPwwIcPqlgz9wFl3KBVLx1WxcS1QiwX381WzzHUtiqcI/gg+XJsYISnX
VVpxGCy5z0xVp9xJjMUfrX+7CEfi7Mp2UNlGCTolWOCDkTTedBT2m6VjydjOUbQtjNNnFA8N9ER6
GpCruO6Xik22fgkdaVLGR+6MjNlNImq8P2Ud68chfA14HdKf/aW9qVkGyGfidXfZs0/TbGiD3dyc
ZcX9oImz2c/F28285PiUs3gO1RRLzEMIJdzNyvBIh7DRjlF9NR6gUC/UCDimViSqxmqzDDQx14kM
zDC1eWSDevIVkZlO3ItPne/G6JGsJYTKIaFsLzNnHP0MzUzemwh0aCad78sDYxgSyBr0Z//La2Zz
lkhQRsKWJ06Rd5wXoDJexc6AGQGG3lECqAj84Dq6iouDPL0H0xifC5LhgXdeQCLxuJELTsbHiG26
UDO5XmZGeMwbfLR9BZbvf0AdZkbAZovAjxSgD+2wAWFbW52TJLW/7nsXipzmdZIP9iCFPfDbIc94
kauxVsOdKO+h2Hr/FDp0DPXdIW6SSybTPx86OYdck5N/LIQHivXkt3EDBb+VETI4Rpc5NrhvHzzg
YLvU4ys32tC2Pck61Mht524tIioyIZC07e3mq6NfH+UwyS6Ujqi7EaYj8Rggp/KmZ3OTIUjxIJNT
4FEPjED6KhGBYo1bfXjgYT6uuXAMZn2UJ8U0gQ5s784zqR9DJJTeguQPR0/hf+EwQBUtdYOIPHXT
7u7G7MqnkcBZ1YreBdFUkcm6ol1L4FGMEZJ03vXQ6GrBZJ8WGtK0uHgXO6Ze/J+ltgPU6zvc4/vh
w60EmKE18uIn+zvetb7l+S5Jfg3g6FJjOyPDxXgM4qZS+dpPsy5XOEZQy136dXmCwMaz9M0hNspt
UDnbyNAp83UTYcV9A8tiNZanlLf/ngObVx2pEFUNiMQ+6pf31D5AUDs23wVlf6SnIFJlzKLRCZ2l
RCz2v/D4ZlOJ38QoWsCFu9pP63X8Co5yvs3/SZ74VpIGWEjmcXfOYt3AZwnY1VKSO3q/jeZGIxeM
1bb6dODnjgQirXiyQMIVerbkw5e06vYhxesBidCVhg971pIv9sDewp0i2TMNmAEwXdhe9O1sw26r
pnxTUu7cTVRvVSQp8YSyja8XKPbgJejRnx4m0QPN/4kLwRz2kZj6kBDHHE6WDKe7URI94osNOtjR
LOHds4OJ1ID8iPrkZd3SlrASeMGIQBXfl7qnlgtCrcXLSb0yRugLA8LP/KuRWKA+Xw5rRrpK6Q8c
7/1DuUDcEM+UHtKPs20scJOlj73tnNmhO1JYehVxt8QWyMqZ5CFS0yXA/gZ2KaR812/Z1lv+ujle
2/jjnsQKE5hPw1UwhZhRMDap105dLtv//jsyq5JI9kq/HvrXzMx91SULPNnzVtiwwPZPnc5qS+dF
XMF9LBiWcSTDVJSqROe9n+Z5u5zj6zibExXJ1eZmce3wlkuI8bfLdRFdM7Vxn19khKdcc3KDupSM
m62xKNE7b1LGaFA1/Yroy1vGEY8J5R7K84SIPTS0ct8GBLMRa6AOJTuj15wBJrynCmx50MlTd5pQ
colFQrahWUfi5LZJ2Mt15hcWow816tdJuQoxL98vmVQiBFoO1TUuJrXIVFSBMUhvYz3Bi2ArgBzM
FyyuHEz+yAHmVA472zr5WiBKTkzSl8e5OgjVd1gLxW07q5uAuPNCsxlb0MxQbxQZaYaFg2lPNXlC
P6NfdX4A4wetLagTN5InGOO10skbRyxVDWk8MT5LASnOeMzjEoaoEEbdBE4F8WhfBgPuaRFBGa5X
rMTWcArPA4EBMImwxf4bF6SLm8lBrlkll36k0jO/J2XQ4TyGBEdOPTCrxznmgLweoA5aAANkgfjC
IER0+J8SeMQcx8a8afpPt/aRUux4+DYsdd9vtQbkLQmtrbMZv4WaU6b4Iejta5Cdi5D9HRXuCaFc
Vut71nl+PjIlgcT3OlVZ9CRvfQmXfxnjhqz2XDYRbdCk+S+PsMsH7hAwWzWIsjzAwpAod5s44pMJ
49jZbIjgynCARHEh/echFZGNa/iDnG8v8EcX9QHRKo7vvCkWts8GtjD/ij7AgjOZc9n/6z3lGwfT
Dry13zurqc0eXe113kpBSnYosGTVTrZMRt2dlirKApNSsa20QKe91UlUvLx5Wa+FGm6vi7tvkcCa
ZC9CYR/OmCjpIKBTlSOMQDn2SRlXNQd9FVRJpJSmK72sKiyVXxER9bPTkE2mMGN6Gyx+2VPkXdKK
KYrMTphqd+O1HD9hQewQgmzHJ8vYB5DgO72g7a2f37A+QQ33n+UU0Lj4pc9nbOOjkTwzrhnSCLQM
6EwKfKU+Xmx4gZD9L4ESH75avTPxsVH8ctIs2pMVnBLgnmxiKHEaoB1f0rWTWnCfBThLtUrQb3PR
CkfuKAsGDNC2O8qulhP8MQci1avdlZPipXlHTITrrkB44xFF5Sf9MUpkeSVrn6zozMnbJCup7dbe
cEbIU8oDeGRuqcnrhsgctanf7Mmu43oC2KYcsZmdRAPZcEr9WjrHgTpF+aDA+LVCyTZ5fwFZx7sg
uyPPaSJrgjaHUZlIsMgRQouZkUIbGuMj55uj42MSLvA3zM1ZICaKUXCfHLAihfYzJ+Q0dZvkmrbO
qHjhv94my+mJoAxJjIlOGRZG18qe82khk6govIrsT/1iDE3XVj5t964lk6YVU58Ce/EWeTibHAiM
9FPEK8ywePnBZoJQ2YR+nb9AoH28x333yDtTDKH8oPl2U/1VJOAHFGiPvQreMfIdtrmaUA5l7Glz
qjqXj+i7OfJg5kHkuSc6hV3jbk/myVDACCYE7Fio7+z0+iTMoAvWfMNDMjOb1W+BhxY69W8l5j2T
zdU1qDII8nS6ZDiIvnlel1jPIDkhyp2SQSWP/zDCjIVMAjKrWvyzsWi2UV6dB7cXxaeTVxaY3yll
PSuzGD3KjIMPjoGHJRi0XO4+I7pIdHmXK/nwG5rr+TBIub3d1NDFJ9rx7V1yWJqYLUNb6TsySHPG
wynMWskB/RD0SYFb/Cch3KY6vbs0Vmk+HSFeVEIVbXBJX0Thf/XXDTJTfaFWfr1GGNHx/1xyaU1o
pUxSaHP8MbpnXiI+nDghlttSyd941BCdHyALNHHI0wMxXK7fgUxvRmgfnQDl4SdtqLNb/QwPRfNb
w8cGz45ZwTHs5Fe3YGkbUX34qaIdfg4Qh+Um4CWEqPGfQv835S/ZkwjPATS2Z9whrNiPXq2qIsKF
EV8NGTrl7xjxzmpT9+x6ruKy2wjZhyChzAqfFr+01eWOt/eF2CT2NEup4HWL0nFIjiSJ6YTkxmEE
AUvjcUKbY5FH7XMysmop1BtBxQL5+6rBEge7CnHJdPawlzwD2sALUnR0v01PpvxI8wGfJfqGMzq/
CsHGe9ONIuT0LBfQiAHndE1261wLTS7TUpvgiaOi57jE8NjAEV7fAK4I5lDIruw/Vb/D6qnk8aqc
Jtq/Bkordx1T73DYael0iSsuTM8fUcaVRD6GXzhu+v30/teZ1RS1fkQImlBp+FjEFkln7zomtB8U
7LOH6Qe+KMDXglq81QK9FqOkIj7Q4NVGEZSpKnY/HqMlWmXNFDx6usKyePioB12snGIxat8xp9+E
G3LibZI7k8Puyaie0FoH/iiqtBx5vCSPkhUYGn9XIacZLbgRH+oqUC3qZ8ePM9WQneUxsNHzrznS
g6znW4CTOtDeYcQAHEoXKM/vzs+bxGnkFdQqPRBqofnVtTZhb76ioE7pfzTq6FsrzX5WEANIwmjg
zTtJG1gsphiHodlld9AYGGsz2SrX/h4ZzWx5IIrNyppHAeZ0pbldiOhYr1EAlxYTX/TLGulXF7mt
YqjnnIZcE5gnTpcg3tDfWh/ye2XmoCDxniHLnWZEmOcPlRkz2lXL24BV0L4UbvDUNCfcbc74KJxG
45GlyYzEyuthihsAJkzu+wEoTvAADlZs4OjYuhHfWY9kmTX9SVZ8DWLJgF+Xty8wsQDasgCWbe4y
vQV5NVTPj22aktLW7u8TPULVuDw5DcRHK3UXlnbsRZ4JlQToouiVCYR7xSM0zXrxCXPLAZYWIYiV
QV+bsDdKOo3rXcVcAPKoI5xeGRLEHLTVG0Skl+KvXq4U4j7Vvp20pJSkNYS8vyFDtiFxIbl9cdfn
q0KmZPyANn7YYn9oRI8W6ty1aOfU5hFGxL1DXk5GyBFXyV3ye5VY6V03nP8TPnzD5gLdJn+v4E2i
9NXJPAKragp3zTHRSMsnVxN4pw9bfDPXu4vP2XxX3WZplTOBxBsSMn+XO2R6UB2nczfY2q0Aazse
JCJJAEBOy3BQ6e9MpSWWf/3JPjeK9h2gnnIB1CssRGfNvoDNW0QerCpx4tj7Edm0zTpnvskznPVz
bXkWNeXOVYJIU49WiGndpb+plP0Wg6nAC7yCbucuM3Vb29oSZNC2BiselqXbROY8kVdAUjz79NJK
SSFbqnFpwu9xR4sBkusEaYrTbTA/3LmAQd4V4p0McP0neGASiqtUlTL8S+zmFZIcPQbGcMnpBW67
iQVSrYXhSu5v0vJqqgltko46hbY7OGqLYXhxz7x5wA6REbwmGc5QXfuA4oWRZEy8qhvVj5wtw+ul
Ja6qOq/v79oyZcVpjS/dFbpDQM54Mxtehj9Jk8ie1RbLO7HwcMKZGNddG/HoPI/TsCZE91dhR/Aj
EsxyZgUFoDXiYdx0c1HPHP0Cv4UUQjAlz23s6iqX892BRhMS4FCZRF9LD5BpvjRQeVuHlw+cw7Nu
dkVxxY6+T2FduUgQImbMoS9CUFiJbR9zHt1R8wxYAiWeqRxARht0z0ZibqQ2VWPdOF5gsFdTV+FA
jOF55Zfm0qf7bsUAzeVL7O1mymkAzptysyNGZGEUNqfntDLxmGHKP4bWq5AhBI5uZARPgG5p/tor
jfofl3+LNE3HQJ8wYsMAWuvBw25s7oH+81pOi/hsz8vuyihA98mttKo9zOoGcZ163XrP2A0HVzIq
ndCpw9RbXxB4oqf9tih/vBckGYcXZd0ZLRauEh9vqtzyDH1MYBWWvqIUvHkHPRrvhm1NHDGDKIqk
6Ym1gF8OBaAc0vLFoYiRtKNsO+MGlQpEmhes6aY+bIlCyh4Te6gN7rimV/M+frs+A/NnZw3mfjZw
E/Y9nf4nm1kkLEslFuJPbmh1z6peMexCX8dT/zsAUFKW6n9KJpyQiITmtQ3Xo0zXMzHj7Uv1k9Df
C0ECdHf4Jrbc0aVyILfV1GhWfykiyvYWNjnZyuXibcmkG1Y7dSC7TRULBVpiY4j2zhj/daCswNvd
nVfeaTTuGu1otdgSx1T3/ignppWSM9qX07Nv9wiwtLYwxsZIuMzRN4eZ0j5qmeBAhRx5oSFM0CmK
tO8DihCU/64hMAuCMDddi+YC31OCTXAhuyuTEr6PpJPnvFrfv8e80XSgcdZVRXUn9FnPvpi6rCQw
AJtVxzYjvJyykDuR5quqA5ebcQpZ1/JIA9WUuyD4b5QaMNZgZ/O3o56+P00V7u+FB2nV9Nqo/hLe
me4qwl2meGRPYk/SrBIZlp+ck5ktg1NEPzkXefoPcbGOIL+IuMOPQMBMfAacHkcavHB5tqnamLIN
IQ4NvxbEUSEp9X2J4eROVtLYb8PftEF/F5x9EsTHdrzecux3hazqtGhxqTH3+zG67tr8mCYY2Km3
6cfHlrvG7Jx9eCjEoLYehWfdmDuwbYMCMIpdMJXNEJkuSJ6+7fBIrDivpXJSJSK7MFagg04fHyat
Khqc2A7Xhn0vGsohfcbLzjL6KRPBZduiqMjClgF6sAyZ3dhbQPgCuVtBVTAgUHru8WecAZZEE8y5
sB+hgrvQ3IBi5ewQDqaxizZjNIJXZTHvBvBMwWN/+wYAH9eRorVRLmCuk4XO4yHmq1lAC6GpWwRN
+Tnc/EKJx0T9aPMOj3C3Sa++uY6/HzhvB6VdoH1azA0lNs2ubG+jo8oWWaQuhE7wP/6TsSmZjhm2
xu6ogRr3vOv8C2iTHhAnt0mPmOV843HWbeVjxqC8EsU+Upbxm5sZrIKJMutFypauwKp2oAYJOy8u
c9r+0EIVCw23WNsimJRc7iIdF6MQnZlfccllFAnD9JEf8KCwWlsrVJuXSja1+OWEaBrfPs/11UzY
piw6WPrnTuYFhRuiOStJg3oiqSbxzCeGGvbnWa6vwOgkPTJJHJrm5P1nX7jsbUB7zbam0XdC5pa/
0WuA+nYtpMNaACKFLRqcBaV/6O7UkOYT1Z03jG2WRorLQwb9Ou7kojpNDVXya3kE1NADCovrQLov
zm+0kxxtXVgNYJDu3YQCvylCX3aeV42wQiTDYsGjmibVsnFIMeZEaBYs4BsIYSgE5qdOBHj45Gzv
q75x+lyq9QPTTRDCbzcysuJRDjr80g8iarvTHmbxOIjo4/8584Axn/ejh4oKRuIiXjvFVAWnL+9b
g1hFJcDtsKSOdN5yOQPAGh/OGRh7adkXQ+tf8uhZklpozFWBJ+wAgCr+jtNYfV6vjZyyyJyFo9TQ
UjVLn1CTxzlMYTPnvc5RdVNDsZX3566K5Rb5Mb64M41L0EoOy9Gvveb7QVJzSo8NYBCFuwG9Fdp2
62MGbk5kfFYcq9Sy4derwEJTHnht/mIagtTMb/miH3zcldksGOnqrie5eZzCI9s8UIHNMP85bHxG
KsdFXcy+zK7A/w5dhFjzFGpr+xZEWmdXBG9A0r/axdloCCvjsJsBj99tjOdPXVI9ijzrnx1Lc1vO
NV63/vvIVKYvVMhWVDEqe7LG4cS+bA6WhE6oiJ4ywCFFth3CHxBNDi8yXmHQEEcDhluNnhkbNY+O
A96lNdmduK1uWXsZF/oRqu7mRT4cbQOeS5r/uDhI9Mu4eS9COmP2jon/+dsaJcQW2Uu+O2b0sTz9
QofwpiBuyxknbtVcHz0EJz46BeU8tBUCvHc9xR6rKB6JgX63vZ8w6NLaMg6RMWNYLe1Q6diwfNW/
0yzUdJph+EOko7uNsqqNyCMKt6/L48rZl9j5njMPfSole4a76jVhguvpDAz7OYKJGuKB+7c+mNoc
kNcwf7mhKxWCrdPRLzeO10ApKKYdSbGZqg8PdVZB9XaoONrTDDKRbLeScioMluEUEkqBOmf9Yt76
eP6+5r0IkBYHxrETFeP6Lr37UQ6mXGtDnQZ1d0cU6u4EHDQUw2HVNewwSM+YMB4XUTjkxfJcdxl+
IL1No+zrfoCR+sS1m8iHidZp+MlOq69GqUzbRrbhWKDssW4BqCjcPjJnZsshWLlGX3whNvuBCd5k
BbZMnB9SzVSqq0cr9bY4GdMQ1GLVzJ990rkgcS4W8vdTBKtUstgrgnDMjFtj3SGS9QOzVfSE11Nv
j+/8OBS0U32pnZ3RNHSpXCF79ZfSz1+ikkTzNWm+a4wIODaAmP74vghboWX7+MT8Utwu7+udDKyO
YnYQf8Xv+twGurY7qaqdDnhlVQFZffXv9SCl9W0aFv3+3YcCRAy/z5wzCA15XjE7sc134DhV7b/o
Hw+UJzXr/bH1P+ullYfny7Ny0KsfR01xAZbiZga6wbU+deTqhJqjN/HqjLthquZjZkbGa6vI2L6e
2Kw4k5GjvCH29Ifse/v3Q73vSfDKkloQie855+YREd7VWcpnOgQjA16NA1pqkMcEvdZzJ7OgDu7j
FzzLPEgO379REf7XGuVDW64yLzFy8f6eImQR0lj2cSA3wihoXbmmCrKwq7Ri/zbj9SK90d5V5L4/
t2BdARENYv5OF/MEgCky14IHe93GbB3NIjFbMixyoQtgkKb2BUFHQQtDcXKja1DlFYntAZPeJibB
v7GxMf/j2/ieclCGdxpaQfyfWTaKUCDEQEu6qMOARKW97sBqhLnaBCF9IHwfnMeY3iYLR5x9C8eY
YEuofVbwc5axeURzO9+fclUxtMujbtCCWga067YX7DSQAiIacQqNCFkF+J0CBjEvNA2NaD8q6AYy
orMFMm/gP5bFmWNS/mzFY/zKhgMgCKd/29iMYOqskNIzQx/eY+Rwea+LvKjAIXH49o0y3ocM8o/d
D+yGQvWPY6wQZhwWNZMJWaamq1gCX2t6cAANpmIy1GHqcqtwy9MWwS67v72nl2yesfmPE6DJwTHk
EuoGi9aMpcOvBRMJwJAfURoAm/mBEXih6E6bX10nO0tAbFvKUrXvL4xi71200MciphC27x55RKaH
M/m5lw2gMRctvFKbHxEeBnMDXfghWTvp+z63azyI1oXsm0/aiGPxJ3n9sTP/GaV2iLftHBf14PAc
CLkVvpZCJ4ay849SHkqAmkQsXTJBzzmipCQ8Feq2qg2UUvgRlgQ/i+qWikhPapXdUIpTvMcELbeX
IfQ04u/5xx5Dsb2P/cuC8hzgvb9Zh+vInKyvyg1Lkh6hJfjwLcK0G1n34NkI8BpaaStHvt8lwCEE
kt25+X3Rip5dT1kBuBMfAckC8CTqS2IQ6PClmxSIuK73sOXVQt56g0j90T9XVoSCYxvvKE53z2wc
pasLDDjAJiXPYZ/ZQPJdwzlMAssStE9QHV2RBAogpX4IPmzfm7sDRTDXuoHZjlaDS/v9vKSQFTwF
jPdSIRU07ATtM3zxR8qIQJtiqoYJp/++5esdw7MazWL+dg6opNpzT3a/kaNzzUF6s2vgNTqdyS3T
REpQmMTD5rgO/rQE0JvAUxrZIBVmhyj/x/pBo/n7BJYzSJYO/wcxGQZGUBUjrjQXiqBBW6Px40Om
q6axAidlB3b0xd/2cKZE+OzUkRhjEaBcDm4XldquVMinBl3YIw/RAThZkWg+qlVFmh1dKVepbHQw
z/NshEkEg7WcIhF205NO0JDiqf/Ue5cpBvzMNxVN4RluV3xwM+d4yV7YBL1rVlKfiLcBGTsk9mpJ
vtTmdGMb5YwLoQm94EsJp7pTORH70KpEyc9DIEHidgpOGyvpZTOy8VfBqFDV2LwZSbH8K3xlUISO
FoA/M6Y9v+eRsJdgVxqfuDxY0fEkdgD7+ReWKEUh1OaxH0zZ4FHYShKZNXsB2nIj/PrYc6+cxbCU
U4jn1DLaacY6MgAkd9C2oMiCBMcbCPHsCXnn6qNfDKcmtRpdJIhUAxSqlwlPnm+Qxs7dhoLc+huD
b2sIBkToRRzVMc01gsF/jyMUs/T9BimYoh19xOiLagGnQJ90kmdG6zjJcQWCSvQ4YpV83ewEFwlO
83lng5mOuI4zIQH94GJ8d9PyvZyT4RiFyDIoZgNYIVFynIO0EUd5QndEj1dJ2rzfp86+fR0/YEpH
veJ+Ojj7pitxbpKL26PEFbIoCUmq34zPsOvdDIMBEHBMLbDoEQ6h6tI5sQzK5Lw/IHzBIDQ0CzYL
8KkpB3Md0c2lIkbFtgRedzMuEpSPUgX8sQgdKw/gc7d/hpWqnNv9X2UvzAyLf948IGmMTrxal2G6
fetWd+go39lGfYNElcWYrSS5oiNY1MKbNhlq7940ecsIG7cZMvgHqDdvDo89ec35yM7W07hl3QLf
Qoc7jMbK3Vu8N/uZoPwZTrgXMzjSv+aoV6KRGlAfGoJkqnoGPfOhO8ziHOc7aMxAcploD5QkBg/u
0ob86HURgORmCgbzMVjegQv5yCYOTmCI3STuNysDArl01QjFsbNRNFphWUZSIbgXPUoymaAhD5MD
TiD9fgnis8zQhWa+ngaCR8WPcsbbo/GNZXdE3I27RJ06U70E9F2Kz/nImfK0dveLjsI8JVmeSBFY
xDp3vWLMKQE/5NVZFVb7ejBKOtywju383Y9evR0BpqPW12iThH3vmctHOsU7z0HOYc92JvkAEVAB
8XtOdrh2UAFL+bJQeAbyHDv982Nc3Tvnfw86jtNVUgt45JtcPPy0zGQ+YIrRxXINwlwddda3vtk4
ZHAgBuuTkD7P7HJ5+edRd3SWYZArnfEFfwkPy/j7xAi0kJVtOy5y64SdKR1ZvBcfs43kTxGttPh7
/h7qtyAhkoTlAtnYG39jr8DiRUiEGEZbZANY+1Ioasyj6SYNXszoQbkvEHI5FHXh4dsIxSs2AndR
yZFWM+4bGzJc6BlhsOmAI94uS5Udi1z7eef/Iy1mQMEvnwBHkSGr9aj3mSa3OI2jiGUghqI91DOI
nARD6iHjjuCIFiwqP9X38xMsql3P2gu5GA57Ng5K1D8IoSOMfu6QxiBRUMu/tJGaD0+Dwr9ilmMZ
UPENNMTQALI9VtI39SafGTJKAAv0N2N+O042W8Ym1xXfHVfU8RRcmENkslHVnujSHU/K/yPaBA4U
nif0ZW37TJIiPRrvYiABc6IFb4sCoKbfMjQYYdGl94DkbpwO3ycUXUVE14NeHxYg//Lj2xPVPm6Z
dEMm68ef1by/RZW4Qe2HpEhviRjRdmRKBlTUEux5pF/LAQYfGn7FitwIhk+RHYyi5XJ6FbiDogDZ
8fYuVsNjob2mlbwcwhGRZMgwNJtDjtKmhrop8ToNcs3Q0RMrlHfTAbEuFUuKGOa+cP5zOSM7JtaB
FsiXnymoVxlt8t2BLZuohjpRJqhMlzoz/gKD4ijn6J06CsyHRj8BTRpkw+Q3/c6bCMxGitaqB4/F
TH6I6dGZS7FKlYQBZ4fat8ZahuLS58NDENzX5BKpeqXTTZGJjA1dTXIYQ/MNxBthmbz5EQ9QBJnQ
d2kOgd+uTQT6s0ro+OPqmNNU5l9CAV7E6Dn4KJ78+S7ibANbIBC3SD8YAoRhPmeoKIlAiv9wpvRI
96VVK2IrVyot2T+lDggWkN0FDfwq5R0Ag4UJ1x+BwOM+DnkV+URWUoCLuawcyDYheHd5tD/M052h
2t5j3lRwe/yTK8n40prqNhkiBy/7emZ/khzbN2e8FDFQ4Y1+8CsfDPUAD1QggXPsUw33Ds075HQo
9Pf+4SnsueyBv8qdK3/yCKANuDWOrYMQm3SfES3eP2IX8E9NSJBjZqkILzo26zJ4P4HI3DfecVDl
x4MvHhNzdJZ3gEM1qEIv8GyGyBBPxXvraH1PlyZ/8Y8R2yjijBlsGfshoDNW/9S635rUXek/EKDj
A/w7VA36OK/lSLkB5yszHX/dfOzBry4pC46sSNKK4ridFFjdlTSbLscsC71pwkj76WatAyHdi0lC
pnjd5zfO6c5uX7l1x8b8YYncxm7Ftxrc9/q9HwCk5RPiCU32uXoBAsQvrO9013H3flDA0eQNb684
p5/vyDAa3pEmC/t/ZC62/lkiomK9wPUCIIvLkp4aQlvdx2fe9qA97tKuYOT0lKLaDgrRRizEmt+P
2U+X5Q6HIPcqGEdB8hEMNuYVT1WYmMlt777gTHnVuHit6Zd/4LAWGXB1Kk6c0+VU3sDu7b2vDqa8
AvDdA9K7SXhgjNhPj2p00oTEKWNErKV59Bk19Hfyiebj63wBReZrd/l/VALDBnWe7D3sBwb1ttCf
xNEXuEfNGW/ze5ubTGKv4loQy4oTATK8QisbyWVbgY5ZG4iLuphLqBT7AfR80F4mW0wFktFF/8GL
4syxfF4h6tpW+KFfeFoXtKZGBVzwLo1SX/Pum3t6EkEkpm9eUac3I9UJ0IIuzGlhbatC6QPwT0cI
08FbFsTVQktrmHgPk8XofGv4j+TE7az2c9jll6VCcW3/XaD83q5PcwNO4QKAapIIfhlGF7DfYYHz
UwEsRy1bnRQquLnjvxCYekz8dZ1Qlizg1j5rxTzKHnv0hlv6MWESKePvemUtiKfKsvOz+j3NNPqm
p9hdDKO8+9uu1qoNWLR7KHhrpkPwdViIjgcwiuGI0mO62m6RoxYZNm5Toof7Fy/0SUyLYHRZqfCy
3Iy/bYFMnCFK7ENSOWH6ubFFnwPFMs0+gSZu+TursAaOLh8bIUjFj3jxOzo0F7jmtHNMjG/A+fnS
/CqZywKoMtQms27r9Pd7T0AD9mPB84BZKagMY9dTIQHIcWXi//4YZGGrBFcGJXkTLX2BoyvTHdPy
akMclaOxo0LqHyDJkxSeEV+hMovCFxEyLO9GsnM8ceLBUJvdV1VOxMCJdp+MXplqkq00j5GgNK1y
947s1L9DkNt/vh0Gcv5lTKFmfIE8Wq/kqE9tBRUtjyH6s/5tmHGEunrGkmBEhakD8vfFxzBB6Mdg
pVSn5lmyTiLU0a30LbF34SML/ntcsjCW97v6EE4RSo34k0gAiM4BCn76eUM0z1JoYNoxPLDjRX0h
CDgrpB4MpVePncfns6matQG4fdQz2k3BByqlqR+nPG5LnqEkO6l3yLw+Aa1YNBrDCoWDigsSerRI
iqzLc0/+MufoZMi3BV+H4Fa7qVWopg/eeWKQHCh6auscdgP/ikeYK2dauWCCq+FepzAv1y3sPYat
Sal2JsWkdduS/d52gXDCr5bNdCHOYz/pxwvV1G3XpvgFAts53HxCYBEJmZ4Z0PmD3fhjSLAcSm5M
nbWV56eQmwiKWh8k5zyFgsKhy8645IMBFOluvSsF9jAbu/nAXzuzJB9G6CRIEwTRWZ52Il2f5Gw+
LnVom3BBOnU31wKq3eAsZxxkd4V3vtwEXbzZBZdDsKFvECHvfTSCs8Wqv5+1tCRoZSxNDp+rKRxj
41sOkvwKyVNr3oxmHgaAVEBjc0Fhy7iYIlBAG2+PLSTSx6rV780YHmEQxnYOtP2iYveCFk4azcI4
R7o6/Ozl4NssBfPL7slS0055HeCMQ/sCu5ulEHNcrOvl6tn35+5d555A2j379eww/2krXadwscjk
ByZHIvZFbQJguU+Djr+175rIXjLa8cEJVm6tEYJ4yWBh5XXgoHfAum/X3gPAMburAWv4HadcxOfY
u2Qm4YdCKa+99MIFDoefkt0+7Gx4PQntGtIiXGN2hnkoqqyWtPLWDMtJmjpcC5iXvWMMgFyjaMch
iqJMpwMhn48NCsa6Zy0kWtLhWHZNvqmtg9Qr8X5wQKGk8Jbt8zdBwIGX5sNV/apSgZanRIOtf3DU
f/fcWm/0NUjTDuzHxJmfwFGzVLZBRfGBDSnOOKJqfTW0rurSoV37cnRVOWedVKwco49di88sXAs4
Fo7l7+tuZxef7LmN9un/Dj5y6W64Xjzv4JPaHvnaHRGc6mXyF72k9uxYqDbjORTIGNd9ewIcVQB/
VYYwvTZin5EulaMbYRlxlJVAfob/w8Cp5aol2kehN+X9Xzxb44w4MZY0usN8/SKYtny0Bv14+4LY
AoO6ZM3zAqM8y9bh/be0jVKz6hdyFsMKarCLeFzAdyI4iVglnUemxENQCrUZfHhHCRrRQqYGK0Jy
yiwQM7aRu0SoUT7r/hl2HeO1Ygx6li3tEbn+tOap+Av3JpsnK3/LGLpwszVv5wGevzTUUfYQbI0J
iqE8pbeO5PTEaRfehQ/tL8VR8IrkWEqutfRA7bcbFh2UvzeZfY0BakVUgAFoYOhOwb/51SGRuAn1
uS8F4FN66TgDKWJ2v61NYTWEUhVuI7C1M+q6mlsRoilSFaEm3FRZpKwcWOyD+4WVak3e3of38UeV
lhzatiEdvEjPcY0lPkTBy9i09ip0IK+PZWcYlVpnIG0CbmLZYb+XdhcVg+m0Uk7e1mGzmwUbFibi
TSUTWwkeYqwZODQTTXed8wU7uS6QeD70rBlUNJ56fuUPkmgH9zlbgI7j0VLNm0qoZjfkYwwkA7qK
Qiob5k/5UOvztCI383p1nJ4Js8DgF+l+V20ii4j8xafl3CbKMNapQZoMq8hCAEtt0cQtXHURT3bm
hLMPist/qyWAB2UrQnHLxqpXdO8z16V//OCji/H2nqMZcAeEmtFEpCwKhMlSOZcoo9HOOAvlR6Ta
yhG9HXlWylOdX6BvnxjOLVJwAuYXR/sygrVwApnvMyu/FLudiBZ/e/zrgWN3igomHnfntZcb/hr0
bvzHjgvPOETj1ES9fuMmz51CCS/JwFDv0ig4xFf/OSOsifXhfkVSTQavTfe4m6dJg5vdpvmvBkM5
157CBctGUrfUP3+cV4zbw6odYiZOw3t0/X/UcMxrS4i7rVI3rZcGKE3ieHjhXp8vA64TTGAfj5gi
dDryJrHsM0FCJLKfcHZj2be7OLyCVC84Jeuci0br81+fXUYv5KIvpUrUkh3nUYLkTa/QIenea+sY
J2IJpqEjDqMHjVFBjJiolU5rH+guM4lLmaTw8EAFv4zKXTlu75kMdMvHyMRM9x1pbKDWiYjBHv+P
tvWOkVKvzPU4h0NyqQy2iwabdfrtrtjlZ5ZHNF6cTXVkutAHAbuwHanVB9H8tqPpCDz5/QJ8IB5E
xBpLlE0kvxL0BMUh3Gf67mN8GLfmgrTjbarjHAlPrQcnZJMjHVYgl4MqO4x+WTpM8Xo2gbXGwspf
dN5ZLwDrg2n2/+QtxQE3uU/FFoVHdL2eGno2QAdpSptGDCyJSYaDEXhJRQdkWc78Pxg83FhXbBtc
9yhqR0SYm3kQZao/WEqbQJtEjv2gKc+S3t0GndwnapIS4sCG4eUGYf59rZRosuF2GD9rvDGVZHmL
12R5CY3SKKR1ZWxIfFDOHrzPvo1/KAMkFQes4/1mAxRnl+kFBPhlBx8QBrvtBxbiusnKQ2wRcq7L
36vb5gRiJ/tkaSThbuoT/3cwxArdBGomE/DtxwdrIHWTjBlJR4fax9KmYibq3zAldBtLe+bPa/R5
IokQ1jTmSMeV4qn7vwuar3zizMkK8aD+QrQoUrVc2H3I0EogpG6/MJV6yZSmVlTS0eNzA44ZmB6r
U/bafLpe4Gv9ZNc+3o+xIJeyyYM2Z98GyFklezZoxvYiRETaWlXJAMWl+tlGUs5k+aAKPVxSB4/R
7f1awR2wlZbezf8DC7tnQUqOKgfOPG7tD01cbBTagAoD8hq1N8e/4LTZckZ/wxb3HKLaOwzUbY/A
sKLFLprgBA2J1CnuITjekRH7glNR5uwLv9ZltfO1hqr0xftNzYTq6GwqUgPdpMkVFQJOkWRAFx+P
14ZlsktwYCt+vIjGoJppaVWt8KtrCpMgA3xu1oblx9Q/Jj60fHIFjM5sLSQhxX6v30SlAr0dK/of
Xj+Jjp4ovMv677/ZA1Tey/Dbp3WkhwDBizDzKNzOXtDcS6icI1uTNjKFGEN0Euqn3EtqQ3VNy3au
BZ9ZfIOaAPovKkq40PuePHqggwGoE/67XdOrK2XxKkJF0RA7sC9t/+qHsB6Z7BNqUK30fjBozFUh
hKmd4AENZFJ4aXulc89YOC60eznZHbGVe2sDAqHI48120gViP6bice/qBFcsyKRMHQhoISl+Xrdt
1aeQoX9+m/w3HaaLQ4IZo455RVg43bHT3ba8N+Rk/c7YU4qAioJX/y8PjFA3POhQRj9DrbsC6W4W
CJmJOsa9KscEIL0AFF+CeLch3XKT44Afu0j654nqb/c/lZ5e/oC46q1mCJO/FFY2HOvuThKGaicO
JLHb3EUwN2ECZhBNF/I2otYGwoCHDVhaC9VPSYL8P8OR+d1nv1RHBzw+AN/I28MgROX2TpVLTpPB
dGxT4SJ9BT37zVk36JKLY9tFIxCA3d7VITzForJ0KAxaH807n5JARtcGVGSGWG4TxSDdi+1uoFkT
xnjh70hY8ciY5RCERAjgIgn9OxcitZjkRDhjU3Gfk7ef/99FUcrl3GLSMsc6NjFf2sUXBnRF7NHO
w4WbQtfS1Qg4VdZG+dB3DKJIIUBAxa3QyuAwyCppfqI4zz4XHsTrmMFMHhJShAk/5OdkXE9/kDd+
XMqzul5gGxOU5rQc9Hbc0JNoRHkKHes3cGQuU+vCKQRXF7cr2MNSaGKPXvSPZFtFr4XPUi3XUzMl
RCw5Brz+XTlvjWNVjfdHudMXC8AIlzkrqcFlkQO1CGWeJeoMukp4fLjx+3/czCF+g6nChonSllm7
+uSf/D5RL/bCfjhrMw5fCh+T7qH6I74Iop8EoVTPENgxQzmOuAsPh5lmnlLarC7qFOgdtxxWxvzW
qlf7FcJJg6h9pCCIdEVcvhM2c1Ss6p8aeuCDbuHrKTWnyEKlfZ1MLIvFFPZrDS735jtUec3wvxsB
95BzsbKb+3LsPeDe/vqOOOrDhwh9QQRo3ouqz33OhBBHJTDS6NTygv/ArrlQm55LdY+IE0s/cjQy
GwmxVL/3UWnX3fPS5A4m2xAMvNLoNKGQBSOHIKBntqkhezW+rRZzFmhIKBEx+I4xls41XyJucNMg
WUjk6hG5OZu8SMRju60HtaH0nNIJ6Ec+sPB3mdtWjr7r4LJZFtQvh+uz3yyv8z5v3YCcLWjNj3PT
umR4u4iw1Ez/jD+4/erQIIfDRhKhQYVHAD0DxoWwFZa6f42gxWPnM5btlSEWsu82aMryheUdp4YT
FL4WPS2Bcpyd0kMz1XcFc5JHHNVybee5ml+83n0/z1+3UV5usuSnW1oK8BMvuAMaRd9NLVhepW/R
zCblOn7GbZBmsYP3Ux9SHyFv1AE+Cz+B3UUVWLNmovdZCrQo9RM1eJr4dDJMks4nIgfdDvjQZo3T
oFjHCp8d8zcVS3wxwuA7Lxwg7fL5rxKOFF3H0LxIclhAO+aYXfuZp68xqtfu6PR02qhHOKqCIBFs
Y1Jz8NmmoQ2iwFp+vDLpl4IDQ6LBP74ykG/BztcTwtTPzSMchG3PBVwsKKkrMh3veT5Z41du4gt+
25FOXtL2R73giGOifX7MUgte3PFyconmDl5PtA/Vnazc9oEDgTNHeYgIjNYEqhp4JTTf43HhLKY5
wRkL98r2XdQ3F+ifGsnRXUBnH81uvEje8Ezp/LO7mYRhWSUN2cTBZBTENxFLz7sGS0R4JyuJbGOw
PXRScsY6MnQvWFxNGE6FRmtsTfIPB9C6QqWuK7+2PZYQvedinUWtAyjZuDlNlsJckF9ySP1Vx5d2
sA8dP0ZLp4Jnwjg3F8EhcKb/udSRiUxH5JTE2y+Dlm5iVe/MebtXFQB+XlwZd9pLKxIX3rBG2rLp
05MDXv/3j84h6Lpz59XE6rr2lQbylM/dfkF0+dwAw9WcJnYNvYcDUxpjYgtza0vBZCVba62CIo1j
3oBjPZtGYtCElEhnvwbC6bv2uCEf0gOOjhhR/1FYycOBlf1WaBWoZ5g07WK3F2qI4JiL2xrFn9xp
rq16hmMy5z4aCI3CKXNHUvkXk82770ruMA3z0FDymhEgZI1c5fqnTaNzfYpCms52tBsmBcEfpvQf
ConwJbFX0VHZChdYN3/ME9lrLtiHmbxgt1xHMNZxBjrnwc78YeVIrYXb+iM5b7Lhz7+7wOSqpwBa
tCgVZEiEgEYAWCVgs4L64Op9JYvlsH9+FT/zIK/Ebfil5zntFEM1G1n90KKNkx+n7+FukSZc4eU0
KrZx4g90s2eGXsL4yZZCaxZRVnkNdZVXKTmLrzMLvv8AePnuzmzRz2UV+HLyYlnSPMYFdyl1siQG
aEGZkhJXQC834iA2mw4EbjueHAR7EfGNAQsTAQbNAXmSwzq7tvfUWgfJpblo0lNjzGaQJpztuT2/
lqdOca7H2w9bZ/WaMYnuWu/zyLvTrfT1HMKT8q+wvvZVPIhejFJ/JtSiZts5y/otlV2IyE+witUj
/Mh55/pFj5Y9a2OFwybQNsyCJ1BrErPtTW38At558HvAK649CnHDqMtHGgyJ0DhzoSQdsgMZcx/4
UPt5ALGB9X3Cb5qwaqsCAClkc6XPbYO7Z+RZ1JixHTefOAJtGRgUBfSORJS8+kb3tsQ7VDi6Dt+T
Czb2Xv6Usps4/ZeHJ4q9MGwmn0g3ZLBOd4ft9RTmdXCVp5PkTZ9q2NATZi9l4kjPFL9LlJISxVUk
lcevaTlBgy9GxQVAsV1cP1OnGvR7VNnZ3x75Zyp95vvcwRpubKCoyoYfZX5PKXlNh+Uef6JYTmSd
Fl9LblhoLhBTXWWfUM4PoSlPNT4OJUEdDbddSBKJilGSxcJMSZjs+mBmtpoEnFgm/oOpjp1MlwSk
FPMOJhQcJadI/PrTojch3HF7pyFDJvwTMZ7OFx82qNtl/fJSkXnCi1DZm+tKwGyIBFSWIeZe/uqo
0hGbzpNfWiagUacXevQrtr8ZoZNzuPKWqWFmOC4ryh1rO7ZE2uZ79xPCk9o4qNq2ePr2r8l14HvN
XO0KH1vNZEpn8zd15hvd1L+xY3DegXTkubT2LB1ZWnVCLde3wLlvrkHB4pc2VbmG69Sp2GA665pU
cuz7iIwB0OZtOw9kHMvtvNQb7ObBexpO/KtpSh1xocXmyK1SHDIOWU4N82kbvI7GmYycK6ybsBWf
Wmcu/SgDP8zT7MSeNtwQZblAC2WzOSYN06FRTsb7MWRRxc+LEaOpjoozbXYJpPg8/w6iEp4S6R1i
btYlqc/VNSW8VNIXlQnMLjpWXoP+YkFzffmPyzuZt50gUu01fUKZJvVKy8EosFoheWyTkkivhsZU
n5YKsXftxsbkB6HwjsWeCWx4W78959QsxnWg0/7Xh/UHEj7aMlZVPYd6FUpCkTZnfOwrq24fSAcv
KthN09VX3tYNB20t7Ii6w2GafpoPnls6Ps0XDaf/8PBT830IitrGbOKUGTJuQIwyKyZijtyNhnkc
z6F0M+coLCo0wdA7/x/7xo7dwSUnRJRcsWRtP6Mz3fP65Vcq3tSJpyWbBImzyFMbLzy7DxZYHl19
zrEkwuQzzOsAkoCGacz+zWwWmmoJCRtnwO7xDGur05jFEMvm7pMa+ocnjfDt/TP67EzOGJNx2A7O
YwvxT4prJxaFJDTb6L7MmRBxghVPFwIRwB2kQL1lnD3pSORwUaGe6I7WIHMXkegkflnsqqvZlA8j
09DctNSStsv7rZ4M5Ku3OdxF2RuFTg+ohzoGcJnzk9Zpl5J1RdZrQCm3HnlQOOIvfZJZ+cIhioyc
XMi6hTyjlsvUzqWyq+p+ZqdaOUBNofgIV5cYUkV0Ek6O0TgMk3XlPXrvaPHGMyYEqMfWXlo0tKcO
t0hl3E7bBlbnKqx9v9HgYCahgCqmSvGkPVqsbMryEFrgeUFmTOu7btuDbzr/fIowUeTAi7SL0IFL
C7S8XNyYrpW1T5sJaCWHbU7Nm2CIbeBNR57EjGQYO442LkgXY7IRa9nLQuZ58ip02SKIeqOaXEgu
/75185clNg913T7PDevXyA5S12s+CbAJqyd3ifuzNllW7UfwhfJ9Sh4Nk1mjGiMPIKrb+BEYdPET
3is/mpZxBKScWn2EUb9p8MSLIEibraCnwRHCC/uep4BZUuMJCuV3I7E/E6RreH4m0uLTztQWfbem
RLafyapAkdM8Rwq3GUJCDoEFQ2Vh2bDW4QQGNdbVVRwokixgFK99cCLVPZfAZJFvTk/DTEyV7MvA
YMVBqWzCYZoW0jwZGRwfANvwr1wQVivEIuH861ZlPRl7wEoFeAaGW3/ziGHFzW6mhWvS5LqRWt1G
ZMHik9xDSBhq0+NnangVdxNvXXvb9Z5MnZ8z8TgXQFkCODTV9ShRv4M+ml+Hb29/VWqNJeIoq4KK
/qd7QPxOJ9kHaJDngJpyWIADrfOTj+A0kZnsLK4IL8tGgS8GVOSAmwVxmsVzD3uQZDMYG8Gq7ax8
sWWnKcd0cp96y0IwXmVseBhD5vY3oIkD4kHple37ShjdH/S07SjWLZa6kZkFMTxHfNGRhwCiT8ML
tn+/mBMUP7Li203eRtmVissTgNKZ4UqGDalDYsN0h3Rt/7qaDn2eWih6CK9qtkRsUtemAk4NqI65
OvGYVY0yRZAjeQ9ZWoTFD9nuu9Nclwi3JH89/ziPgM88BWUajICB+8EWscm3VMi4othzCwS1rbCi
PnJwYaiI6z7gQqyyyoyhO7x4ZfIGXwXoMD5cNKX0oqf+l6ukssi4YFlyWepQ8+VDMTafPqT+DYxN
xhvh+qCqnKRAfEW8HwxvvRs0KigzjzoDke7t3tgvY0mMEnCxyA8EnLjDuiaw8/Vi9PTKJlOqH/9j
UiSU8Lh3rTgw7DvPT2kmRcfdbrPgOovDFhOWq24UioDRYUjSVIfZIV/wN1jUB1ffmuGluzVl6J9f
C/5Va4L8tMxBfxUOkWUr1sS3MlH0mUDhKSk/QK67tw1lyRHZtD0VMHoPYI1R75OH7h4oLzcRyk2E
U/Ej1y+yOOWDFpGjS4F/7JFSi9bZQbhpK82RM5neRdQ9UQGj527a/IaibNVcBtDOo4fUBVWGfi8B
LG6ZmfFgCFSgeCJeMd/emhF6IWkDitFrU4up/gQszcp/PXTXeO/L4fyIgMOXNTbsfsM2QRcAhmRz
eepSMKn1og0S3ke5YEEo3qrwZ4clGq2uvPr1ZBPPZr0yw8LG1vuXWNwSZesjvfxVrLxjrno4aKVa
iAyv9OuqyOf7dkzbawuDuXWTiMCZqyO1xyQS0Ls/x44FWfQth4qfWLRK6zTuxyLIoOQtrTLKtxk6
Nhd4AX/9/QL3EhNAtBgFoTGYxKzJfVv/2dxi/yzzu8+D+FbVyFZvdMamgDaQdRoTdITu47XK0Qi0
6MgYdOrKw/FWpJwDGgSJ1C8fE2xv5pFFU7ZBjOITqt7flc1ckFKQRugxqe8XxBJEFTtFdbRvcZ4W
bWBPslxgt1UBiDi+fBXRzleU1R68y3DP6t5w9d1BLh0qkUiC/7jpPndnZw0Rp+NzcnZYpUB0+iTR
BzrBUL+mEZ+/CSh8BgrK0aXpZrMCWZ3RA1APesqSaC1ntQSkviVuqIgS802IeslSx090RMMm2DSe
OXmr208JCB9udDw+GwYrmtE+lCxJpzPMwz+++x0Jh7ShPqPq9n/a1IaI3PvemNhD5hUv3B4nFMwN
aQYdzdgCG2MR55g5xalSUAijFGPSgXgY/uhroQWxHsWolJCalEC+dfItwNBjfE5PjJ6g7XYZ7xa0
BERgiTHRKB1LDh1S15FIG2iWPO9mKjJGSTMpOzG+rE17eAj/pnZF+uKyI1So84MomcCKbpHwi/6D
5IwowsdPHnUt9iX2CBomE3COiK9zw5Kktr/QjIlb4V3cISTeYoYOmtN5jbOKJAP+9QxTEYxQbTaC
HBkel/x2AJ6kyKhvs9IB4tZt/Ap5rgVefVMPgdn/s7+U3UmRF3Ga+x4O7dYgsL+PUqPGoG2qN8aJ
RZ1bpCzNln3gdRcTRUb0+GJADCQgvPVnqCqHnjRRXqhzsZODoWLQwvzgv71culwYUV8rT3UYj3Vz
l6eOQyGzf+hTBCXvLDnZNsog1EO0Uj/4PLmEJsyv5kVgmDvUP93xkUIBNGogFGN5nMBEMPwa9e9J
I5RokSEtN1PZQ2JKeZWxxdzWT5mdiYdOQnU9RWFP9TdvPIvC6enbxJ75Y7/JW+J3/eqUSI8XiSgx
Do8d5xyzMhdkRGINhfQiuc9xFKJ7wkmEi9J3UM7obDSp3fkb3EcETP1w+eC9VsgVt5MrjR6bT4pE
6VnR7q0HF//s2h7om+raJH2eoNO8G5tM2wfPo0UBtoLGBa9Kb8cXi/rTNZYnVLz+HRi/UyLABrNZ
nlLjQY/wioKE8IzTS9AzeT8aWZTe1UnyTMRC/c9Y6bDHnTHrmJFxzhx1YQqNXsNSPaTFb+xUVUp7
uGgkRJI4F37OdH2m6c3DbpjiBvnYXBQvW/0S1TE6OVEGGFpAjL/OPk729bBaEkrwgneQ3moFPWa6
590AP8+D0yIlpvCoiG5VG9TXVzwevPtRyP2yKOG1HDtQOKzaVaWVut4stihh+elbL6AKDwhyhhC6
PmtCGfnMO20RaW1WHTv1lAr7KC8uZfdGig8TnM8S4dWvU5rQuLSKOv2beTiTYaB1G330gGScHoDj
yHoho37rnQFtkEQ4dnmoK7bwSlGaJziYWDn7CeHzZYTuRek/NPY4JxPFpTERVISqP8xZWhQLI1G1
HhDQfc32eZqj5JwLJbmR9HaJ9dNTTBbTfYZmQAwV6EeqAQVzvHiv/5GneZ87aR/P/LkqnMWI4QrO
uXZndsY4xOqGUPAORwIKaEFD4rkdfk9/mXDuwbDKim8Xm0xzrTO96K+UFFahVCW5yq0jFMLbGeWg
bne3YGfUh5X5zwrybEkoVj9HTMC+TTe8moFFbOkbEPDCGYSivgXcOWE50pSLh67uD1JWCubfN6+b
GJfBwhxZJsEhfHqu9xfFTHm/wsJZWGf5J2WMZ687cVUfvh8op/gvYYjvSL5nP7F7T7qjSggLEcBm
MBXMmWnJZjNyxEX9cPrCRqgFe5nf5JzSaSHWLyjNglxzrIowusv5ugbAzrksw0Z9SpON+zo7b4r9
9JvSRBcHP80kQeylr49VRjx2waDESjgv2ZuWHoyocWQ4yWYuu933LKgOTluX28/UP2FO3kEGSLHZ
5zptrIreldDoV+mEqUL0pZqp6NmeMzGoR9vwBLYYDPfGQw49+sCZONA6PIChicgkKN/nwFumP3JU
wVBn8LugjPCY3XNB3qTJamfQqEMdEHOiL4mIo6GkEiLdSNYTzFbdL6q5tCJptBBeCsEMRmWuHV0m
LfemhZUlcv9Njh5Ey0QlwwfkmiBTBsP8+ickVZzoxf6JnZLEvFCr6xj8m9mex4EhowN1iEgD8onK
NN0WJ9GD808/T66rXlnkFMMVgFIFBUvbSehB+AjhwgF8JrH7Twx5tLBlW//8cAk3jJKpdUhpVk4w
+t/ct/4DiQP1YrweL1hFElKZvcw+vLq6J8+ag0V6xGtqp+7mzMQ39I+wAIt/8XutxCWf+hFT1zqU
Ka8qDgvimt7fsSDXV7CN84EoaWXgytwyoIpMz7mHMQMeWPkYgHfqnPr9EUH3+thw/ojjiRG8b8FX
bDjv99MjcH7nGRKvpAkb0G02msnEY9+qxO3fQxBazwB4E4GXhTC0ProPPOwko8xYJ2d4JB3Bq/yw
dEeN8FLls2WupCoiEknOVoyshXolaA5hEhJPsiz2gtSP1x4cKQakuMov8nT9k86Tb3PiyTiXx7Ok
P/TQS7IP2KrMgeQXeYqWVCltSLfd/bGse7TtfeJ8+Oz+e9GDp/yam8hgbISmqKG5PCFzfDUSVkPL
N+kVCT3S+DUoX1wyGMY4ZceJjHRkwF0jAPcgpSzzO1LtGb0h/28pIIciX4Q9emjQbv+K8nMhqPcn
kqk8qxdcs+5mL4x5UWJ1/YftP6LhEZBJZWzQ9+MycESW5G/L9oxqeHKoKk+gXRtP+xI2Pg0rzMj2
LXJUwm0frprDN/xSXzD0dQnl7jfZ4U18D/sBReLPPXjsnqhwK5Q242nbNzS6G+GvbPAVsUm5INrY
l8Wb94JQTASwnsxrgiGEUYSusd1MhJWmTK1OtIMfifpRBoN7e5HHbtLIU1Z+cWtT9c17ADCiWdHN
igDr4WWJue4n3D0FLfzsAGe31hxbK0tLK6AJsncV1OV9+FfD/C0tLsI2KH7G2UdZZkJlYDJEMZe1
Ogdd+37bWXTwcB5NoVv0F8zPSs0UcTk9wjR5SuwE4FTQjzC9jmSNsulFDjfnYO0fn1U1OT1j/yTC
9A8tQSaNE4nEvWxP9B7ZTVe9Nnfht0MAoUtG7965Wx0KronT3WeYvk5YezbGtCRhC7ONKPtmrdW0
4xVfxj2IeWo6H41nMWGpf50eIl7UqInOSwXOefWitGdxG5ZCiybeOJm6iifCZxPchVg01NL3Q8jh
f+hyRHW5gBlHyRvtBWKzfVn6dcMbPPG088oJUfgS/72aRjKGjbTaLQYGy1secRmA3B32LMFmZqU9
Ba+R3cMR7L+6oIlUssLJpCHUq1I8idDyHukFMDGLfi4tmKZC+1MzYI3G9z/nAQF+8v3hc3zy45Vx
pBd8zI+yJKa7vmVg/HDm6BG20xTGlIjr/wwdIO5Ir6HkoD4zI+FdAbe/4188t5/zNWnKwBjCQQBc
mjYM9Rp65onythrEKcfAhxTBYbcZYvulOHe8wmtz/+e3sjrKaNXXrPP/Wc8nWaiGQld5li6Qjp8X
82bypuUdHK4IIjWfli6bWXZ85DJKQtyyGqhOr1LlIpaZEoHk5YfqXCS+vSs2fG3X/6fOp8jZHsyr
h10Zvhv6t/mNcWHfMKDkUU8nUh6+QEAlsAHkt1YDc2g1R0yKF5vTkFzm/hsErc8W1mu5utGfEaeH
0VXA0gF41SpdEN/37kb23/iBGmlbsly6rbcZ89rn+HgGLqXIk53B4AlrQ3+SFa49//v4EzSr/iki
rxBLc6E0a2+Ee+BhoVRBwjERiDB0rdmBBitwsE21q7oZ620nlRhNLqEeS35Amy5cUw9RTPJPfQSy
Qt7y2Q5EpHa0Z6UAZjsubqZ4P95gylr4PF8xSI646C0+UYQ5NMCFR5t4fgF5tC/EC5V9Pvo1F/EE
LxvwCwHrgoM8AqpS0FJ6ZHPWk8B6ASw1aof633MmxuaK8QyxqC0uOzXGFiVJvLm+tdnW4tP4NVXd
mNHrrsWswDvuyKZl3e7dk/WP5IMkWYyDIqfn+VLzJNcFY63YLy9wMJDSTQSutcZM1bxBkYL/6G/m
e5niUFl+KjHjVtbptFqaeEyGJJXXeEnSQLgLa9D7kQbU/ASxnXkwtUlOoaThvxp8/a4QDkJBZ+DQ
a+7OG0oOahg5spUIxu29I6cj/4m3qnA7fL84tG5rd1PAtRHkCAODsABWyIk2NI8TA+m/42EmU/CV
72374Ok1gH3NY8ZOKt1eqR9bwrOsG8rbOLH13/TFjlyz2c1s29HB7K72toyko0xZPKEA6se9/2Vq
7Q8nmHrpDwmfrSkUBzBIH1dozF+TEPMbbH/Hxeg5nyxoa+AAfKTLWkx3ejANbsOarQvmhzAYsPKb
tkYR/mrJEyM+bhJYIi0K5C4jFbW9ok+LRLgrKFHXaGPO+csRpl84W91BN7jrr/cRTuve0mDMqRA4
fhiyFWUK+V4xuKCWxniNgvOh3AzJxsc1vheBmTKKWh96SEZfnVKIP4YwP4prtPnGIqp5Yfb08ZKe
7X6ek6EW5ficMfoQyXYE5vI1/rW4t7qxfEGLsKT/DfGR/1r/ktICzNGROm87+Y1kU4qfW05kjMTM
tj9vmeGCBum7qYvqvp9cBqO+cgsA+l9mOcTghPIwDQs0r141f96jPceJ2iQdiTMSPReR9RF8nA7Z
DLnANBzhHXbKmQb6yBHlmbFify5bH0KGWOAMch7pwPYXPuHqJWPJGq0ezUX+eV/KkBPDFxsclvQ/
g7lX/rBdzLUDHez/AYRiRZZPh2EQshs7MGdNmnWMF41ku1jE2ywPSrwLYuQ17w35zggDuibePd5t
ZJPEVd7RVsQ0MpwNNc1u4p3kg4QAFN0YYxe1tVpSN6zBsuFQxeaOwiV4fuWP4YKl75veNAKA4wxv
JgFg0vG4cHMeGja7WWu5N3zuZNDhYnR8P8F41YAplDev1u8MVqZD5ZicGMGkTFFnZ7lhltNp27Hd
z35WhCGe4Mb8XBXQa1Dk2rrgyD4ukedPngoEPwriCXuAVOsfadSYIDZMbBRzz8wEctzQCdy5YSp/
qMSVSlklL534QUG9U4o7wRA0HTBC4ro1xCNzePVvvaDDfTdi/r6BI/qbx4ctpQK77bdMqaHZnR6q
o2AB47s7FYzhZLP6Tv/8YMwLy7qRPmIsmxpKi7mhe64Q0mYy5AHsXPRbICr9O31WzO1AkwfMZEnw
f6AL8/QkLdAQz8l/Fm0DMGVfg39DLLV61CkIwQNr3Ma+cXi3H2BRnokzB934vm7qvvtFx659nJa0
F7lTqiBLJe2uh4Eu05nEFECMZf5pPQf56sp2I/GXay9KXZyqG5nJ0vGTGgctuo5wH6WWKGDpoyIY
Z5iMQrN+4qC7YC2lSB4wxkKwzgly4Smv7ET5mO9+UvK6FOmWiI2jFepS1zMUr00LnEmUQtQ+i9NM
y6tUwKAXiioZ9gRb8efqHJkWA92MFc0hTeyEWYDnj8dTuZ7NQN1Tiw7Jfh7NGIh4o3aowzI8hK3H
9XzpEVn7JTraxd4chS3bxymQdQKWgDXk2/0z1jZvLJZger9QqAaQ3H5LSH3lZxx3empRiabVmw/D
abuf1uxbrSUnidl+buVOZA58z06gFW9P4Zun0VaMqk6HX2kUmiOVJlwoNTlX8rEDu7yUhaitWaaA
bpxWTAaPAeHxhfXbCd272uV1FzIM6YDXqBhmYjzzu3aBPYHW7rgNlmaYA6VUX5H2+4Sm6dMTc0Qt
v/BNi/pdTneGzZPhce/wz7TfUDP8HYsv7UqKKSMqGTEzn4FFtPJYJdjBeGdwKJ5UErqEKoXQtYFJ
jIlwrGC83/UtWYNlRZK++o3ZMD+aLFDD/KKdDCUKjrc+ii7C9qzldVJ4is7kMx1MDxN9RnNUXUOS
v4tIbmYlooZs7mETrXFiZp6L+uL/KZN1ueUZcmEHEAEGjS644Wi2jkVV5X1ffjysjNWd9XTQ8Lqw
tiltfIKL/NB61XyAUEph5K6cRMzLtpiK2wCh5zptMDk0Nw5IJS+Qm7+L42h+gZHMACCcVIVVpYF/
mWT1bCUn6VSEnJbC0LSgRP9fEBIkrOffjYKLOstC7N4m3IehXOQV8y6guZJNnknLkv7vTatyTGL8
mcxSkAXuBx0l5M5XpjkIQawe6GvmqnjKxBHng1S7GpgWTtIKsi3yrsq08KLL2MSGBQMZ71DhKsS7
di9abuZztS4nU1Xp+BSB9GYijqh4WD3XCSGjFSzh3xM6cCnv5Mes+19m9ovb8q4nNqC9ETszLK0X
MUYU52q5uR8536xZvpQuI7P+uSuysmNOorrypPkjl/2eaWnLjETSqlMOcG2xMkuDdSC53CtmbY3j
827SqCv7wPz0rCs9CvcPQNoJiuJw71/8J0oJBnqFYPLAw9KPPI+y6HpTcFrP3uvU+i1hpnJ2keR8
bunslHbdSaIVdiFwk25ESFNbKpzFUvKYYETH3mFzyMmB4tboMo8udm+CDx9g+qZ3Twlpad5Vnbtx
D3wBupXR9Q1KkxdcUnNJiRmJ48K5vNmUdUR/Nag9X7QIyZkQ7HC5yNkLstN5vcvTM1lsN8kxjSUU
6GT+cKhhWBlfb4YOEA1EJ6hDME2PgI76cAa/Gxt2OmraMu3u/VTAfIFjFDWhFMRXXZi6Xzt4Rl2z
7MqH+1EyFD9aPjq7/rY1dMF1xfdUVdnukguM7XhxVDQbXWAHjSzYkQNIp+/dLPr07sn6fOVhSPyw
dRO86eHFFjpeJQg54tP2xQEkvg2kFZIJWwc3c37Qo6Bm1kYkLRQcZIBnwO268SNKVjYi9VLpF7ou
ERzixpwJ18hxXJ7zljq7g8MTUtYE7Rz8FVdOMTFzJ2xgBSM0i3q/9nNdfqIaTDh5XFZ3zE61Q9/P
28kbGnICuNMS1Tp2DnY6y+Muuot4wgDRqrqYwFaebrU0QF56YRsHLqXSOzGlxwJaa1ddC3rAq+b6
x8JsHYEXxyudCYha9NnJtKoJ0h2leu/LPkI0motNFc6M3c6S17khLtOkUCV6e5fsCUjFAL6+7xFf
mGUId7JoqdZ2uNTA7XEGUk3RnJx63NSbq3SQWRq0/HNSpIjRZgDJ+oc1Oq67VxXATdRjq1T1ZEwJ
0HMrB51wD81HjogK3hEc+PzIi0sxEK0Ccf4R9QXKIm/s9Oa9XQ0UWeJM6pTlglcqOH80bZKKxdj9
WTWty+xbs92PaZlcIzJW8ZBCVNOg0KAoS+9FyCVWYN7kxsDHpyKEnZ2gYY1cpWx0CooByi6+vMeR
Ysl0hn4XkaD3rUIySJ3IbzoUGMYwjCZZka2zAXnmxvykxa3bjdl8oPn2QMgdHLOJMl7QKh51WbR9
/akUbDnbpJ1/zdceSW9Ecr8Bw4d23CqqqyoMDaWP11gws49Cb66pY2ew36k4tIXgXq1Dcn3qIoyt
Fl/MhdHW7r1hXER6D3rC+yf8nbNRjR463N4wkn3MHCCD/ErgNcGHOy84v7IOWtG1JHhLZiNwrWrs
LtU9esAsfugiQbqSKuM8inZPb70XTz/+BlPTF8I2YTVR5KMKF6HQQvYTd8YQK2KiQ9wNcy4VY0P/
5ZS+lOg+uQNb8Tb9Ix+49o30I/bxiap9DJcjXaUcQVwZiZdwf8XFNBETTvC8Cu6Dz/aY+WWo8Z0B
dQJ8HR1iAwXijz5A5PeLUJx93FkxUXSUPbv5vAQ1ZrGZmsFD+Twzl+9tdjTcekaDL5mMH5LbzFzy
wU7Z6dQRuKdm4mjSlvBUh3bDagFM8zVi43xAYUL9m1VrNZ5diqxwEkoNTHer9WDRua7w/EuqITLo
8bqMRMWlplwkGj6qoDjYMMincGezNT4KY7VVuHmzB4tr26VCX3zufTghkzY9toBGurajmfjjGNAN
nOuSUIlbm2dRZYBq4+cWEQj4L/BQM+QzIdUOckFLy2AZ+2qZCh1gVyEUiHgQhioJeBBOfQl4mBCK
Ix1/qK3Kc5ITAc+iA7fbkMv3wJEfYtFmjdtYJ0KwGdd7wC8wYkjt2RtZVAW3YoxEbWfG1Ycz7jZH
XxIZg1Ozqimt+aLwUuw6v6j439RAIB5voKIxsHUSjGCVsFyk0MetZeNPUfpdyxj2EbIcfvhoGpJg
kQXIMt0MfU/V9NNVwj9Z2SIr/KPlsfX9gk8PHjdTSd55MlGWgUqeL/O1K67ZSEYJ5DPC/4KcmUYk
TcePwymE8W+0CnxCNseCImLRq0am36ReCNb1y2UgUojOXZhPW2DyFozVBPWoT16Gz+dIsNrE0ph4
k4LJNQiZPiUcFY2i5VUe/d3y9/C9OchHOmX2bJBv1icEzB99uNmkLICDdM2tv/bjMOrYY8Wt4LCI
6OzxqOD353jBR4/WU4gqBkkgZLNpuKMTJYmnPTYeYwoP0Xr3vz4gOR7gDnOTdx9pREsmBhXIfrnO
IGzsaw0Uxxd5Xkos/znEVsN7j+qS0z/e9+Wv/sM+6E2XLODBZSqn0H0WoyUUYapYmXK9iJo/d0/7
iQGZbP2zfXeb7meZ0EDu1xFePQw34oNxuwgSEiRyPB84W9fwaIZeakIGHm8sTeRyyBH3FInFU434
QxItBkVIMAh/nvD50w24xKp/PIgNqewyo9RsujVFHYXMGl4KeIFrDftN/SNRHRZFOtvPAujhw4gU
Y7IsbhIyJNHiu/4UjoVAPtgmerwo54Na1FOVnrRzi971bneLlTJRxXwAx2NXOdGVPFUWy7jfbRjd
EZEqq8ipRs5QF9F2AgmaHkFMh1Q9lyVGni1k1CiUDKMzod4S/E66WGQ/5HZ4Z73ucnZJSzYbHwV+
mRSLi8S2tRqBNdGqfjUe3O3CCqJdSzmjGvAdNeEY+lKD2QiD3yqk5aVhZegKh73/Bo2zwjDKf7tp
MCOnzZVd9rLsbcejkNuaLUimYpHCk3+a9cSu1y6d4SdCLJkaeTCGZs8lvamJRQfd5zpTaT9xrJCC
oXT5IXg6L3+JYuKEmBkPlfkJa4nwTpRuyY15IN/Y9dugJktzcHbfnvz7GPenLnJOYx3gsvslSQFB
MbFgDUbbCzazs+7eYgsOmDuklNFQN56Gh4SNGfPjs9NyatI7cpFt340f0/bMY7WpQtXry49BLD+k
Cgg9ZovHx6IGwbDB/JCm4aSV8rPujzBI/ILdY6k1yr3hMDKrr8xVein+Zi52eS0uKK7GxMmycAHu
EWhl4TpHnU2MHebw3Yut+IZI4JWWZzj/mjLgJ+wOtDx+QQq/2Ks6Vzg5Cma7NXVrOx2N/xlWIqn9
dN8VV27cTJjnX80jcvCc6HJDcsoEqZRFOE6QhESj6AFazLoGohlKSo9ubhkEqKDSHJOOfhGxtI0T
DBDG5tawWLJeu/S0GRk4ELnsKlApQx1ZvKOANrIXFMGG+hS78qIvFfVf3ZqLvFXkIf3AGuTFArdU
xbTA4SckX71XG/Hl//6p8ygARFt2iNP0JJoVh0Z9vyCqlQbmI5pCwL6VS9vdq9jsDwiZj/fxz9nt
lfW64NF5SgTodgIYQHMobNnq90jueyYdksbWfYKutfaYB4aEQf4if21UWripY0lOY4IVVqv8kNcT
9+HJhoGsmMR47T7oAF3kD9pbRgUyl6dqHziWPzY18p8tBfFeL5x+2c04ZMwPka5gxRNU75ofq+lJ
ihyeV6vH4q6AWznfUQWjYsKT42Vb7MChuLcSNefEG8XyhTrLuhcQaweXXqojtsIaFdzMkMyjLpJp
cDV8L01JQoixyjCSdOfH5/uvkV6mIEeOL/5rt6CdNhuSg2YAJI5wRqfhx84JE2UCaY2SfcLXKGI8
SIGYebkKWFK0PAg7nco0I1+H9CBMUjCmXLU8CI9aDJ1ZSnI3BIN5+Rz/gIyw7nFuAEES9qb2M+MG
jVszUwN0gLy72+TTzKljZh6XYPi7B1k0p6qIJtE24fUZ+jbMlvI3BGHHBCE8r+qmdXMp3OMMP13v
8xsxpbY85mE266y0VA8kF+kOJxPGPdEkbTzGLqqYqsqodzMM7cMUERCGot+5m4Dva3BSBpqWO9iz
/HZsoSvAcW57k9VBZtE1aeTFZqEOG5Zwb54bLXeUrTVW+b3r1uvJQ7Ikoc41UCG6mv02B6Rtme4Q
UKV6Kofd2HpYQHlEwDuv6wWfqYqitAazVnYyY1iy7Bv0YzF3otsDCdzlfjSWF/CLbbvG9cJ+nXWL
jFYNYkmvNCyKJT3C2fe5BNIoJLAXia3QfQFFTXtz9SberN/uptOiR6MRAI9GPcWCG5AQbj6S0Gmj
Gfdr0gWQEH1SFoPz5qJKgbbQbRpAwtFQtPVwEbYRd96rhGGI0Pjca/LjaH/ncsSUQqzHIsZJfe4R
XBHy5hyRHRI5lvIwr7Bttl8tPLJrRNzzrmUIug3uvBL41EobwkQde5KDKjL4dK4wLqSt3x2MOGiS
pGcRqYs/C3qZBb02AoqfPLG1cDdYSfrGS8+sVRp/IEC2VkoI/T0BIDn6VbnUhh35dRuRJ9EDj3kr
uePj1TZomDledYqc7YJguBZxw+tbwbYkYaPsh2O1wD8USzSxqkPn3IPZDVL2nJOfQVR0RCIRuKSM
K96VcDo2ObfFHV5vB4lI0cn8BR7WK2DDATuMIOlaW/K7fIevaCYI5w3i9d4OBk5QfGsfi40mVyGi
WPcSEIBqie++e5u02KQw2oq/5IQsPUe8ZKtXsISOoObEl9qp42Wjp4DJV3UJnZGzlSZBgvf9ucfG
la7jVg+bq6aBdWLjiL5LNwHp7/2YjgkINWones4Lcx7Mo4R71FtGTa721kmF3Fd+t/utuMQtxBSL
awxtRGyVCwCczAnCpg+KinQh2F7U1/sOFTBEIew4v8Kb/Lhi11sUt6jbJwFbQjc9hOXz3mjyD5TH
cTNm9aZ55fcFLKFECRw5QxYKuz3i79Wks5iUhPjiTSTEcVWH6GZfGwyTvH9XP07Kmk8fHpqrSGOj
O2uMf1qFXSvNMZPKUWEjRmkYpkuDFy/S33XWVBZTani4KmX7CYwY4kdn7FEI/uh7nEvoDBeAm7Oo
dDNBxd+moQ+m31KTm/5B9AguGcTcsjnNEo1tb1nN7ay9DkKXI9lu0AxyS78mDWQOWjsJL4C+awnc
/PcPtmg/q/x9uRm8qMgSDZWl5YsxFy1dqw0FC2vQ7f7NpG4jiGhV8YbY8mvAxpjabg3S3j8v4Q9h
Eco6NKqyJ29jU84Rja90XxWJxnXXtmYMqfHlL5z4RE9y2mbie6KH5CsIDvsP7Zw5TsHIcrOQgLQb
QsOrSWzY/FT+5XnTwfDaoY7vBmeV4IODe3Fc6C2p7dvbYvFDurc6llZvyrRAVpqvGXwxSgQ4y5y6
GSmaCc7sKCpu+0w5IF+biAELndhFco70IaLiIhJ58wCacwUC1ggww5pSO4RbmQnUP116hIeHKjKS
zBagCZR08lhKeGUzX9PVCVpqetMfzx2WTWsdIRG+fRoz8ncuj5wZRjnCzzubN6X539WhPlsxoR59
PneePKWdVswtSNTrFGCexGq1smlyYk1/fj5gEK6K2ZNoLVDSmQ+V51Hn5iQyUIuBSC7nyWJJCBU6
cfkpmmVCl3RvWW7nynQovTV+Zugc2iwL8yyuq3XM2wg8zdbZpcJULeBz/R9vo71NU+l6DNRWkseU
RA5ZWdk6IaKRnTFk7dJwBvjLEHc7WQ4kI7d1yIDUx+3bP4s3kSYtLylaq56QeCnrKRE/EP7w10n/
qICj8o0xz575fTjd7dDjgv4k4H0mamQtVOLxnm9Zx1+RlX2psWO1M/KqEsVd5nlzF5+KhAZRl1zV
8XGWTojSuUHGMTKqFqMiGEYMVjNUEyaVb7PzGeBb8+c4b82EcGKf4D05EkjKCOyLTMF8/uzdWAPv
PGYVFpF7yzd7cGYtxV0ygc//cnsJJh3/eHYT+JZzcg/+uS44TjWlXxGtTVwDbCexYkiZeJGDJpVZ
nM8MU7BwHtXBiRh/hB9S9CP38DlwQj0Q51PIWq+Vce5NhwuqT1V3CWJYA/VFOicu8VgLSUMX6dZt
ZRi6fdYBUzCPJfCoNb0E1DdVpVc9NOOq65SKYLdXUr23XWeOU9gMhaxOJZGsI+dJIuJqz+HWjfIf
xxmwdCgLp+WS1yCTt30AGWdXNvGILGXKFYp6MMiLNGGy9c+UGmxmgMX6gcBZbF2rN739OlneaYSN
3VfifEipp4qxrX+5QYE/B69++/O84w7AV2zu6qxENMDG87gXv8dV61n7kK/WFZzu5XRwRwoK011e
Nz0hsoZzu3YGY4ccKng7JsXgYI56/5yBr4hJJsdIM1Wj1Pr7WunR3BOcTg0sHi5OYrTVnHtqi7H2
LJIfT5QaayxzDt9mI091/UksYoDp7zZv2m5UPBE7c15ephkXnbpKpUruFG0+jCaze7Sq0UK9qSNe
xNKlWw2seIxZF7vtJGXtStgA/NYzZDzylXeEzpL/+s9B+EbUJJJ0kZjbrhbNBTbSZBjCRMs+Bv1I
/IHAAAyrTglVqs1F2fsCyjczYD+yFnJ+e4AiqyCgdAJnOpGMWxlWjnJPj9nbHps/DZNV6prgtGuf
0lCdXbBBVbKwOlB0aW7yErLccn13rhChqdNpiyT11qifbRMrVxM2npyV/ccp2w0aCQfuscGdmlt+
OqUVpgrQvWxZJ0hV/VTqJAe7wxwmiknlvAjgkngECMD/2tXoXUFMNW7IjI4bgYxDwKWOMmSuHQA/
dMNNlHRNWNyRDbD6x86rXsbLJw0mZ/yzUrq30tzjD17jogGtSGknq1mKvkQp4gPQl7fOxD4vdjZE
IUcxHv+wtZpowEn/41LLrjj914IB9RJ/9GUbLx8lVpbnElMAnJonUO8W4FWN9Z2L6XKt4UacBkbB
wnVMrNzhQvhSJzYpZ3FB4V1lylQlgrVdEHcsNARR+bRjMuQR1s6nk7jJDghJnsfkqJitJDl3uVm7
rCySctYwuGEtDInflpVY+0srIQySEL0nIB5lDcYSy+o2Es56nSUHhPPWuNC5Wep4e0F2GGqC2LID
idhR0vFpE8OD+Zm9ahAFWgt4CLoiaq+BUr+YkjKEkTUhRBfKaT4pe8jE1iyDUsGjsrOj3E0IY8ws
cXTWUt5gJ0gA947/lH4UXUK5wY9pxrKWkl+pQ0Zj6QOMf9m72OPs6MbI2gn9y2zMbLmxnAryOsEn
AHVSG5Gdj2lgay9Up7nBDEX3H0ZtksJ2C29APpQdoyZb41iTyhbJFyLbdwpE6fueZTtkrMWsjkEG
+6DNn2/wvGy7dTxScxfXcTw0QbtUNyY+nAlejaunvl25KQ2tfevuzi45rgxsPWb9fQql34Bzrph2
k6vwwnVppVM4NdKwZAb0lMIIg7dSlqhiqdWMzHEJc/gQD11wPF5CzSwJE4tTRmfYrdoPR72dPd6Y
460nvaWd/ZA4FyUt4dx1WO0cgy15KfUET07oZESmJnsHhjaRes+3kY1EY3y92xZZRKWwVv9vPPr6
yZ9JQjsdksvjolYVriAWKmPltADagLv0oUoTwfd5CsFxVfPELOqTy7xef3PqG1dGnFsgp5NXOOcY
bHlNSIHEA7Y5Ni5BJR+MM1VxyP+MJUDVQQwBukRj4/CzwxKGfghaepCPT8Qtc/+PXRzcu6uGdWDU
haT2GL7SW889jicj+zJT0UxV7KCtCTbuJo6P3O1inFsuWBdxgiXxwyhRQBpHIoZsZ1Zk/SE6Mvxs
xucvBoGlLIw9+sR5ZOy09HOzfocQgAVVoctvqYMB/iSpxBCk5P6HW5Vu67UPrM1H0B28//C5Ou+S
qMLc1U2tb9r828x89yW5UYYoJVzW031Xn1mt8islm9tergvFSWC3fgQ27vZCRStk6BW9qtu7NZ2v
uuHSGTEhTX4A97jZWzhb5QVF7FKmZJZEWAHE9NR4tLFbwoLtwov3566LdirZx0UIZMG7sQJMUcAw
fGO1sS63MbEjNiA8Z7rv1pQukS0G2EI7XMQWPe83F3Gj5CBWgRVfHiU5hbXq6btAFQhz8JlRphGa
ooj2fKqI/jLQPCKG8xH0mlkA100myerdYyXXxGAoBjm745vzmAHGm6lK3ytHx1VN8K7OxZAnzeI6
P3M2hswcirh3A5jm87XKYFwrHFmglQLopa8R8OulQqgATB3V86/ajwJDwMLRjpkeGFcVw0pGmq5M
e+cuJua0i6Ejx/OY/LWmuUc1XvXhwqRvIezuJ1JzTFKno/gzj8heE4ay8SW90rbMrd3DQkAV5cOT
UZFB4+rhNAqTRHmv/QFpm9R7H+ZT1owV4Qtufkc7Ts4b+8q2UGCSMD+eFC0NOzDpH4+nu2Ru3d40
7OQOojOH8+ocjV+3YDvxPj+oDYvpQ1q6XIjGSm0WUxL6IQsUO5ttiDlHYHle+GY8UVY1edwt2akG
L5OxeHh7I8j346lg4O64HnHJo/dG75DZMHc8J3B2L5HHIIJmzfdXPSPgOOpp3FurDP0ulwzj3UFQ
2L7Yc7WsrnhW0XfxOGBrA33FNASm/MxKpRj+E+lh9vrR/R3nZ0Ky1bgsml4lRTi6XVh7VNMf4A3L
79nHW3sI6NZzZLvWwoA2daCoNFG8UUrPYqVECm6/OojYm8sCE4j2xGPM2CecJfHJVSi8cbAl8I3Q
aFGucxgpiBSBTes9YZwV1sIAHOG42vlOaVELScnrhO8GFooO/eDvwfFwMjOkzOfdT2O6FMpTASpj
e4As9//09hncoBZ8Z61fXYAd3+zvAq6/weKwjiQd4RqKY50EhBSnIWLy2ddAi6xG9N/bRkAzRhyA
pU0WqvyPzZHlW/z+iGceGVyHsS4WmQPH5RYoVv7zODHJTovi9CVR7mjF/PAkiDPWvxSR77o+kohr
qTsc7G+RwXvGE2/d7OsFAE0luzkQqKYYTKGyOnrnVr2JqE+kFAFt+iWuxbr4eH4LpNKg5GOl7djc
Ii4yGF1oepipouTmnB/YP3sn7T00bmkqI+GhgzpKqbNoYpMLHcB6/Zlcf2PziXWnx1mXdHH0yGjD
zp7iOT69PMK6ZzeEJxmTbwyn1xHbkTHTb8Wh3hlPq6+Oq5q0VutxSO7ZNYI2ilsYR97EEFl2WR5L
DAADxJS+d8Uf2/eCSogWng8GlTTRlXfsIBsPsS4johowzWHkIS8sSu6HS2sd0vAJPQsBUTn3qoY0
pm1pum+63e8JXvzwc76nG1+rI6otWn65Gx/iQqp/WefsC6KvoosoW0+PFvhMYYeHCr5/fvbeCybz
WEKwvhILCSaIr5NvBFliZDfJtwXWZYgUsk0fqvx7QUBSsBDKflj4+H3b1EVekViYIGkwd/D4P7g3
OEJ1oeEDS07WdnpiefN1sXr81JY6Q9Qc3DXnxlx01JOrgmPbqzrd9RAxsEPZiHovtNyseQ6Goq6y
A+vz0NpKP+1O1Ms4QEKWsr5yz3Bvk1aL1gwBmCMMFCQYJeEvICwgFQ4Nf9uloGecmIKDP0plcXfK
Zwud3x3GxdVyy7yBZysgDLAR1ohy7r9kesMM+0OKDo5UkVfH/m7uM+s8ekY4jLaGS2gpoNXpDxZl
VKPDPjIDDGndu+aRhsfBsjwf4jWxkFG+GxZikpPATdbUd2DDQS9TwaWpZZnpyMoFPJ6K3H+XIwLo
CHDwI+l8w6Ri8k3/uQiTh/ADXahoxBZBY/eqfc67VFEdamoXGYGeyHiuwH/GPK+poOJ85HWrE4zl
m5I6tiWVXov2bMHhO8eHP80ZqBHsW+fYF0te73wNBalg2bblhRJ4h52Hv4aaIzUEq2JkQ8rglqm1
ncE3iEC1j5/Ydnxz7CdKnG8+Vb4EE026ks0SpiQQC5NKt8JBvTcUV3crsQ3qL2a9Beokfljl0WFS
V/WCU1b3etZi0a/4OTRlVxYUoBsFffcfansVo0fBlbPaRzAhvHG7ToAiSUVxUIVPBjNBG3l1WxZy
0M7nvZVNeI+rqQjNWheDNSNrBVfs701YSCrxVvln+CVjKFJefK1gl70rTbD7gAkCYGpsu7AvhPav
511ynFjcTuKeHH8YI7FURUMa0JUlczkg9iZ3PCNJ7XPvoXD9Dy1z5iWWKHoJsN3HwRDr/LqNu4N0
za055lQKwzZJLleJwryiDjN04S4GQ0WZw9+BeA5+vezAwQzVkqupstKSxUtfeGDDsebFJ+g3SbeU
RWqG+2oM4m0ItfotyGNyyHZOKuWpCbjKJpip6tgmxMgBl92gULDFVHQnnXqUSfoa2gVm9Rez3dtt
XtSovr5ndIKBnCpP6tNwQD6FBXIJ4Q3gxJAcEVWBM0JbmAQRsbQbDMm+/rGDdgay/q5/rzcf9/tE
QA0t3gL6/Dg9IsY1ZUQIVp5OiLdTPvdSdnHBwStRqgQCfztNiSOdycdBzHC30RkGNEOnKVaqYBWF
mKhCvPVVJlHkOtxyeamNvvlhOhzt4vQx+rPRpa6i31pqU8jf8Pt9Ad6UIXns794yJkeuGMMnULvs
/GEhHaEvmV2WpK6zsQXcH7Y9+eG6ANaZgAYgtL75PhndnKa+o0S3d72ExhK+4642WlXu2tE5/JGU
mYQ9r1U1D3sOK50sCJja3hJkWyWCF5uewBdFdhHruPo7WblhuMdV0tDKXO9EB/+656HeCvAgp+/N
lfjr5XiC9eB+Le6CtDmQ5MYYZ/efDxNzstmLrnUNXAD0PWd6NN2QumoAYuHfR3eQw/b/xxq4G6at
OXa9+RUaNtJjZQtHg+tR//UqekZSUM8sd4actJLS78x865vzE0greHzUa/hsqrTLWjok078tNRtr
foq467/i5aWjCAyUqLTegFTtwvOoWUf+KMfOLL35nI+z9+IJFBlCVYXDMVr+wdOMI588iYXJ/Wum
9IUJKbsNkTJQP+7Srgo8fxRdvVxAXSdYmPdtW2biRuFu8iOHnrMNOjqoz/Y2fKilwwRmYD7Ezfae
1l9ZxXIvB/sOSVGWFrxo8w6ak+iZHq+I+KBTtuSY4koEGF2yz/128PgXhYVdpXejAFv82W4SQrLT
Ck7MzkXq5SzkFiVzy4nRPuibWxnWLuCQL9iW/vDYPQZDtfaKxYrpXfIWPWBZ0fAFNLf/Cq/dAYRY
dXxiciBYwZLl1bOlSo2958lfCX+r6X2k99pLdJ1FCY/XkqXbJ8ZY70fah4N98+5+UGbZj7WJxfPG
g/6ivTOOS/lQgwxY3Y1lMCZOukdqkSw/GoNijxEqO01DHqLIuJ51PXWuxa4K1qsHoLUMVU+oN5tn
cuYzpT1d/HJMvQ33OGKKwII8rudGck9ZKqSPkASlhO1vq7DofmNtzjuSIO89qkUa0EezJ1VhNIi7
cX2ZeGF33kss8MtsvUXkzgQ/cOrAHX/n7w58S3NuJMDRS/jelnLfI+M/o6rOTGM8x/HuBMQu3S96
qfwPdmXkRzVHD9zpKvjmlcetL/HX5k12CyMA3nHs2HQ3KQdSx1GumDPr15uaMyWI1FkLTmNXsfkP
0ZVQi5+GYE5f3w3cdSxM04VXoM2sArQFKMOiR8Xu925Hp6Id1ocDSscrudPc1p6QFCAzVfTHvnxu
eSBUCVNe4/Yy2I1BsDjDw2RZLOt6c0luIjPe6UJEs33iHPn3qPawyD80/I6Ow7/MxFTciV8zLmy/
aEpQWoKwE9q1P4LBEytL7xBy1JNXau5TIYaMTF6BZA1dGbp9qhPMXO83Np7EhSxVIdy6JSyi2Y8m
AedeWFy2U5BhzyEnBVgFpfmkJFOwifixHI3JCkPEyEqsr22PMyUxS3SmjGjvRKljyY7+e3IXFBkD
CsrafJhk6Fk3VNUsqVR+3CZpw+nxSYZ06PCTR6owWLWOZBL722HYphIQe+BBfFncn4/rixmcbejR
0VVLLykwcrkFyz+ONUPf85dTjCKYgGzNVVIQObUBjejnThOTQSR4AaqYs3DRvjS14c+uXr3C7j++
030VCR196+8U1DGMZejIzflkeyia5lDIZmnhnkKcbXgP40NVOKNb29jX5eLiJ197NZeJCgTYKOs7
+ljZwGSgexy0xLC5tzXjq2LlUyOSop3tFg9B5A4wl35PrtxVFzNGtv5sy0+8KYSZWP8GyyIQRP+0
56zYzXIpfOVGqQRfAe3CTZTk6VJfzH/qESfDsA9rzsiYjbCsfGQH+DslOXD6qGRL/JjZIr3G4T1V
89QX1Ef5u4lESIHbVliF7kKzbGTqcJxrIfjRypSWp/3bFMIaGCVreS3QhxsQOKH787z6ec75AI5Z
Cabyb/VOY2bB4JSMBxTjlXohtZMb7/5v+wRV48WPKQLpJa2fUnm8+yVbtVBB0VCx8wB2IYvUQVI+
l6J8g99dcT+VaN76pP3lIg8b9wqtHHZ+cNORCdazErFAFy0o1XFxDiHORF4iXosmB8vTbmT+ljuM
LfKF/L5Fbkm0Mpnmapf7OCXp+FU1N7dL3P8KPK3jDzkhI9szf1HJ2GjSsVE1eezURTDD4OwUEe/C
J9fiYM1t/j3FBAXwnhyOMajB8CjEyRFXxWBR3kURZG/X7Mkbae1NeJanWmsAId2kn4ibuexWeX9v
g/8yE6VYsWN/snVFGU1opMleHJwMgV7StZ0OH8LeJw8tUDq6nRPVQjFC+A/BNglYReBv8EjsYdrp
TVkzS44n8QA+6JrPGtNLZuEQfPkIEovkukR1HTkgZ0qbOMGdrRlCTFrpzK4Gyjr02IBOEEMfT042
reUeyX7D7KJJUTN8LwZxIX1LaNGZxrGCa+E45v4KNt51FEOaihWxEfM4TJw3WYou8cHMV2vegnjd
cichXh/edez+LurghvLh0Il5xm+Kg6IxqddjuTDPDWN5uQ51PffOZMCWYdc82vs8VvywHP0erUX5
L0yneR1hiaXhRu5YneP96TJQZ9O86f007OgyUbMyMYVntXQ/UW8Do6zDtUUJdtbp5fKK77I/MMZY
dJAbDbjZsg+PZzVqtazl8r7W8N2vs4PG5jqtyiKLu8M2IYYiHW+eR8mwRC+WYcQiC+gNwLRpMOQY
EVX1DvN6cAbisHOBMSKxM7cXGoxnMxVKvAfI/+p6L1fcRRuBCzBcLhyt/qy6k92s6/df1rvYlwxp
OL5ywhtMZ8EQbywahwNkQ54DQIFvviJDvSxfuBMnk/+CZvcIi9p2Tl4kzvA474seOsQhi7GX7reX
5Q5XI9te9ojafY3D0E4uhlUSKg2ADwz6T1riXH//5yZDm4WKk6Ryp4JwaI+3meQG8ZMQ9xGgeauV
7KUyQkeSOIK11Yk6tjNunSLnCRGv5d8ltulrG+T+CMfWY7H7NNVUIPIjNgRL4LWV6AYmB4PFCUog
8qXbs1zLVaaAzmxoqTyNoflsOWyn/LzvrwKeTW+6/+xyq+20TR73Ko/SQqVazQ3kS5K1uZj8Kg6O
hDGoK+OGNppIfGYLdUTkTATIIxFA6JseXO9HZDdydTnCXOxoSItcTRbjUUp7chbTqhi08+RzcyIb
RxMH46ZkZPx80mcP4n6DtAYEhud1lpT+VFqBMlQP66/rbbS4PTJGsrhTAssErmBAaT/eXWXG9W/V
VuGuDud/bYTEDvGudYw8EFzrFD0GfcogChrJCPQ/g3iRgkQTJIYgb0WAyVt9P9TF3wM00uyhWJqx
J1ifC2UnsVwi5K299IaHavE95A1FHk/2F3rF8sCvoCHwfw3LjHYsmJ/6ETEYzpkfte1XwFYIXYaT
OkuLroJNrICArWsvdB8fSgbntINi21lLFN/1DfikTF3gin947Ds3utpP2X+PZ/oC6S9JVeu7bsDE
siq3XGlafHjwKeJaYVUIXs0HvklO122UGnaQSr90Js1cpsgeKsakPICEiVTwJP6CkUjUCpXwWxW6
2uolEObFY9XFgHNHq6cPbxZzgxNW6Gg+DyNFn6FVsAGMSxJdC4CKPuGpS7RbJeNmQEXwstLDGRK4
kRAGeOHSJAhdteFk21xLicpYWTmvYtQb/eRKxHdVBc3NyWbFdUyzQeW0oEr/WsG59o/euiiiekuV
+ncevdOJ0oHcCk/ZgVx0mmDUEYBJ1dZROc+FCi4Ctyfv6+uglFZXFuLzaRfR89TMh/6rp59avcqi
ynzO1sso/6hqnCWj9UVFTqcdW2vgKckHNIy6f/xE+3mcALSHdJYTKYAmbrURbhOXb/5E6JbHloDZ
GKGn4aWaUnUz5+9KjnC/cIcmCtPFtgoHg6MhFh+0Me+5O2ExY/Wl2jfICWiHoLMNv3YgE9BLarUq
zJqOMXzQxv8dSaKklvyQ8UMZ7Y+o0JLgfyu1dM4XJNXo5hK8VKLxiLCiq3Pkw/z4B/EThmU/KWIv
3a/lKHbHn52X9dhrX9zsc5aVMd0UZykN7dRmS7bSQoWOCA74Dvyl3ilZLK/x+eD8wbj1DHTSuyrq
vB+6eRmJiFYxEDg9SO7MNTkkgItaviVWTgOCXhKTvqfiTevEgxHlAskheUImubq3Osc8uTTsONI1
2DGDuCBQQLRfKYSPdvFUh/e0tb1HTpFcC+T/nYYZ6Si4QUqMxlI6OBNe/6PfO3Sb4OYOhlJy+Xcn
sWMd6U+1XQROfTpuCWflOYodrBJYLwp3DjXZuwG0SiC9f6oX0KlgjlwMmr0mrB8TRtVO1vKpIq7p
TEU52hHIz8Km0/CgI3DKzDeLc4ZkMbU0R6PDw6qcphf0ktyPf4fPiDMJGMzpf65bfCCuET3N/rQp
HjHmVTVhWnGoyNcucpApdUeQ+jWGsfwJZCqFXst8lpjj0hCubcuxUBf665ml+t94ecmgu4+lQmWa
z+kypaLPOIyWDwt/lj6bat9kENEwqIId9T9R3+b69XEFjVaDlpaLIlmqGpl/buwbj1Kw2Enl2F+p
wsO0qs/OOKPVLsmEFgwaZIDYZ6oro6tjCAfc1VXENjn+3ngkDc0CkWoF1Kzz68vQg7x5yMpAYZ11
5JV8wZMiekZRQGxWC4sjO5McUYdhkcOszdPqW4gFDdAzC/ohmIBHNFc7fNHZy65Z+U/A3SyCyVV7
SedI66gwyVWvVf6qgTVyfZC4uoyI6GT1ccYmp+GgJ9ryz5MZu2WYS7FA3HFL6Ofu8l5B7PwRDpQw
pVO9rcYFJdFDuTrC4fZYYUhwJPed+9q2xYgxVxEgimMjfKr3PPOFz45NYqTsmLZYNLftFyjsEtyP
tc7MRXf6DAqYBf0C/p9xiB52UWmpsmvVvKxKNO5TTKc5K1jffkWNiHRJlpzAtFDUzLoFwWPauMCh
ze7upwtTp578ch9LQzX3aCXzyowcjuBXBUBqZT5+MtnNZ4keUzgVp3D58yRbDXXFyWmzrnLzdZIM
i2K/FIxX+H1sluU7UV73YU08r6JHDqDfUs9Eqa7MV/flscI41QSu/PnhZuQhfzw3Smf2BE5mAPCC
LY2+UzmhrRrvfhRkWoVs131qGbn4xkFvDl8eskk3m70cJN6bAf6obIn2a6+5SAzlJel/XzK/Gkom
yrNqPpPlOMGwE9snjukO4gs0ZSxmfDz1m7Hv1CGX2FMa5OTFXQtMb5P7DambyZ7U1hysBvLKm6Bl
V/j3WS/FAxmWfgTccHLw369V1uQiLcpefm8khIGq2wNFrv02dtibhpL9wBLMHKOZp2h2akWSr2b6
yqGtFCOZ45GEfUDrq5F0od43sdFKavzvXKYnNZZDK+YkJYs3CuxEVe/dxcbyzFH88ev7n4tirejn
/KGuHCeqBxEjqDxIRAMAI1V+ZT9sbOANSgSogAUcxo5kJ2OdkOA40B2csgH5v4pkxcHvQwSk900r
p8jsPSILjatALMPruswEpV7EciCiHNxLHMsmKxHvlRg9eak4YLn/ggeSluvYQ5f/e5tPT1BbtzRW
76CD1Jn4wob6KYNNTz9S+PtuAtBuQR4Y2RqDdFPFuO0R0TfG+zsD5uxaop6s7xuAnTKGiiDkPx63
sNaHnZIk3WQjwpJiKI1Tcmui1Ugj1yR2MKTatObJcObwRa/m32f4l4X2lbGnNC4AIXxj0jnuILgo
j8jR696U0e4o8zENLHE1MUgdhtRVhW3/scvB4ZgcEBnoXsoMdpOMKtBztyO52ofWIO80A570ZB9w
ActlSAkf0CN30q9Bi6KSOk5I3DkSAPj3oV2/ridq8FxvJNhtc4guTYsY6W7OM+J6V5ZC1bQpqCas
ca5viEb6bFHYVlOCkarQwsrQn8GvPjSn7KJS1/IsyJnHC3/9jt77N3GIk/HKbgLQfq7hfZtRgM02
7RVZ2iCfRlXWEPW4YlrZX7A9aWIMejNpEylr4GnZqo17uqlLSOXpG8B+1P83Uv6orj391ke9XAQS
ocYXYTJqP8ooTfTdxIz90f6Fol4XLleMbVnbqQJ3Ptb+jjLegRm1AiMjitNvdLQlAbWdEX8u2mRJ
BEPzfmfioFsOC2CWCKK0/TTdzcx2Kli8rVHuRfNQw0nm1fIxqBHY87ZqrrVLl7a17wNmChnvQjJE
65j3sEQ2+tkkqkDUnx6Fw3Rw3DjP0PgMlLhJVJPqPCmlGbRLHEddV029YtQy+DMSa2v0V13xE/hr
SrxvV4KWN35nURQ1L62F8RdwyMumZZvH1smrj/Y90pj+nNQkOFpi2NqTJtwD/AbbgY40uTOZqZF7
f6GzQERKJ0AYPREulL1DfGRVnejftaZntXp1gbPyJ47UGSxU66nqeuJ7LeF3RQQ6NC9nmdZSH4Ff
X6V62fsUrSQtnQiJIcXlThrj8vyNrPzF7N99joPzu+qYi4koDmzv60QhYH0B4SHVQpC0S4zLvSjB
cITP0Ynop3/iWWHbKfrt2W5vXxc2i/HJFboA8xgeZ2AmcUNEMSrzOmiDc5t51LPA6hPKyOF8Aqpo
fkOcBtS0+UtmNQ4JMOg7mg08IWoQETLfYUVq321MwYTpT46sYfB08bu6C+DtYanxzc5Ts/Kj/3Kt
6EbSS/DJJE2oO8mPS/FvDTDWAT9gXsDfrC7sAewb6FKvkAWAyAfOdqFFmGrhfS1ZANhrRRSmP1XL
QASOEQC//u3eipeKIbBxBbGAp/wb9ttqKwySBzXeLI0cY15v4WaT75nuaCWea5hfM/ZZv5IPuZd7
amwx5RjJ6r1cM3bvUTSi97U3lsrhwuMyQN9u4ti+9xqWsf1FYJcZcTkQoyVVaZR42Y7hQxY1X61Q
GGB/1KCvFwfeKrCgTmeMw6BujrNA1AnUcnMeNRPE/xi3e3yYuVO3BZ4AfEwUhEO5l6M+hFpXnd/R
WoebOONXS5B7M1WdTsfTpby6yIrwiTqCXzdDXsuGrgaMwIPqT8odn9U6Vh9Ae9k/spJ5sxPYtfx7
yEhFfKYu87d9XgDHfLFTd9mfXZqx4gR1up8U+As1WPF1Hd25cHxWeRwiVxCaYqlW58NANP9L4BQ+
hYoqpou0jzZFEuV5LXh4PdTz85uhj0kHfTtWuU14MA/jnIzJzZijRiueQv1wQoBat4QrrtjNNXQ4
8e3s8tI7KKCscWMDxtolMZRqAOmGnvhbEGCYQPWcbzsIkOWoQ3ljvYP3Ry+woAWCWGdiew1qSVRW
c4iny7XgMQxzLR8py9XhJVZycyIV9IzC1X2BszwzJwz+KjrvLzuiOFM2he2JkpfEhRHkgLuDXTGF
A9mzDN877jEAPdIxZui/mypgvVyr7lAwPdoafy2CLAVfYoECz21wMbsu084wZu4O8oT1qXAwMbgj
6vytP1dKduwmTXThaMgHlAZXEv5QuM71wLsmIih9vbbgmVI/QQmL8h7cKl2MXAs+znaEa72F3N+w
37iJTPJad1b293AJTv8rkSZ9P0SAmQRw31NxYmdV9Uxnga9PC8fVyOqR7S+d8a7BKr7+NpTZ+yIt
PDtSjvuTC1VDXTKJFMS/CSJEl+gjLzHnhIsVz2yJBHpB219sON/YV3VOzvguF56CKUXTKgsodNyb
ZeV2dLSxormJO3Qu5BJcWTGsaSq1hkaumw4Qq8GtpGoJZVbrnRmy46dZZ/5LT6h05yPZVzbDeHuw
WA2i5h2QgKQv8e9ZZs8apOusT6sfVCvTXMu7I6O2w7iYEVc9xLes0sxlNIsZTO3Nz5M70ny7qoYK
1OBU9YI7aT1CgDHiWOLwsEN/2f9Y8/mwgtFID3boeZjdOwSdtd5ro59SnBO3t6HmAMU0K6URs98G
JEC354/s7LlcWegpLB5KVkUugKLAO9QWEpLqPJle+MtL9ntPuFj2fEp4W77mTx+TompZ5iPxePtG
c1nBSxxhs5CwvxUlStBjgH81VnYaVX2zod2fFAK9WmXZ062v3xVLj5mgXccOLeZB2CaAXqNvhM/f
uX6EKZ9JQAG+i3EMLwPt2MG+klv24cxkFS0yYo/6Ihm/T71zcVlFSBNugZBVUUQ9sN950SzL2c8f
aN1ANDUhihRtHCl0g7tm05Y79fLfg06xmiO89YtVLNNKGQ1rPhpLMmF3xK/8XOAWA+HpRP613Kbv
H0BgQmEV+Ys83RDLAXTmyxe7qLO/q73x295hJd4HP4GxBjIUyY6LAmLBWJj6VyXyyowzqZgSKp5u
BSL0gT8Z0qqFgefbWh6UjQMq/C0SZ7dxJcu1n96gougnz5SCkJ1hs8Z01+4TzDvnSc7cvXIJHhXv
NECcUdNjtg2OfKmCARleI12ZjgEF7WMpWrkqMFTZ2nyEuko7EVb99pGfsfAp51b2tNou1Ha+MnII
JZ8vAuyThC4BdZpvlsLNkgf6GLK+g4Ho98cw47nNgHKDaUfwRqjsgmrH/QIZnU85ARnr9uSJQGwC
AFrTFo5tnj6pvCOpJqD8dkACOzU19FPd8UE/4APpqRWUqBB5TzXsBca+faYug2wEuSk3X39vJtZQ
/A3oAMq+vHKTfmC2TrCN+GBo78ai1jbw5X92xHqMMZ3u3nSdHZTB9rZkY0Zia8/8fFaEmBKz3sP8
9MwVVkXOeEir62eEYTxRrUuXSKVQGcBoojIlZum2RblfROANvret5o9xv+EfOvxpgqTtJfBpx7nT
wDoxyc+tQPvEZaE8sxuc9hejxvkbDTcGriSOK9wCTSRRM+cUqPS4Di69AYPc8FCt/QQ2pVUcEfxz
bEvZ7fJ3Y1TJ+i39oMoKxURGbnGHI/bTxiMivkIoc6UXc1EHshYIRIOt7miE+HPBHbplg4NCRo+R
PbaStd0CnTfOwSd2Qx57Ru44fLcEZpaWPLWKHuIsepfcF4218l9u2zcPBB4ZSPD6Sad68y+wYDwo
PIlYW/pUIt0Fxn4LMHO0WdmecRdc+x9nUHGnTT+thUFOLG2Z2moefZ+cg+3ilatsEqOwjO6/DENP
eH12bDGuO5g+OR5VNy+kle2XAjWLo1/fCPPV3MacOluxp8pFJ/CRnySQ6EUiP+w5IXkT2SlV4GuY
ZpuK7Of7pnEaM/53mbyKJnytW+5UvS3Iji7kzJI3FhpWZRQ5aHmQTF41geQxSGLggWp2nO2CP4LL
zBJ6Cq3xeFXe1daAzuyp1TGSTiB5WpH27AJY2xm5gDdt4JEqHSosqbQJ3FXgIKnRIIA8/EAN7992
EzZQBRWs+Q3AgR6o0gqeHYlMY0zeNm+eI7eGHcB0Dl6Hzyth2G4/cCvovFIHI3XguCPpKds4Lsla
tOZz6B8XG8vzKdO1UBKlTny3OHyF2kBUy3Ahr3FC20qCba4KUtcldq2UGqVjahw+1ctkMGM1EVXZ
QlDbDaGeWptjLgPU4Mp48gbs89TAmTA1RqTGiwHF5NKOGvzyeelF8OrujrEeHe4NPGywoQ6cnh5y
lhEMYLFuWw4ItcpGgQQClHlXPWCdAjCB8qg6Df30RgNMP08bztGrJQr4vlghuovILYIcs1oFy/5R
I62UoS7Fj5eWzur3wsG6cG2N3orT1o0Bv5ZDTUWNEMTCkWHl4XVeInstki4n8w/SCpBkltQzHplx
ETvAsyQOjoTK01T6HzJB3+tZt58ixijzqfdgjPGtMTwgRCjWlwGZeZzW97HU99ASSxxk7Fa1iSCd
m0c/peUoZ7vs5CpmSzTHue+Qzn/0XDMsw2G4J+xIMonrSPH72a6mVeZbcykuOtmsNr8G+2C9fOIs
rZh8yFNXkaNEWJ4aK7n/bzXRHCv9SVBOK3sCY1AJOUF9SUrm4nk5jXVFw56a630SeAdK4dyyYXua
6tpB/rK5/6np8Hl+rp3ovTV6iCKv5l/ncpA48uPWyQg1uoMRnPAqmR/AIl++k4PGV36D30HVzEqD
mxn+TF3VqJxseENhmJlPkq1UqqmgmjrxZfVUH6JbhlCaDlafsljlyGaw3WlQLrSZ5dE9RL4Fhhcu
LDyBrCFCXwFm1Oj+uHzYJExanemf2UPs1IhuoKHODOIeDklUCj4dGavC+7JM97HebvauV3vyVh4S
rpZmJaPIfqyphRZ/nazjHZXE5q3IxJyg2qy5zhmEVJHX+Q0+l6ug5GtbLCfY7j/QNy6s3Gox/Wjb
YzuDNXGMz6DK77dB96qHSLJE6Bd4qauanmI16qQ2ZOSETpQPPsz9wkwGZ8E5moZqvaNHY9u9Hm9R
12gzoJqrT9tOsK2Kr7W59f5L4S4NMgsmd3TTMb1vv8cpfj3OT2PJ0GzOd914oV68rYthhv1OUNqI
mZVQO6aXuUjHDpi+wqY0la4RaBlCmalfLR0oEP5PtTFIuUJYFwVI1ZSZDeCRB1/gi6ba7hc/q55D
wwWpA2ApG0U8uwNPmRnPKpuzYbTNAFjPBsH/WRulccNEQnc58Iw2yubqRrj1cBKhjrdWmjFepT6e
j+JXUs6vfNJXtgLWXKBiSVQBdSO31ZXHnYtoLjhk03gsUtb/UtlOQQjYFVg7Al6JM5HbUqYLlCKD
SQgj4o6T0RHYDwE9v5QbmCdynhJYsVoOCgRjRk+3iTuo1uarxZaktdIgPwLFHpkHrO8NwqqzMKwp
m23MNIZMSuXVKrEV3nrEyJShyb7VJe+eBzTB4oyBKiM/wAVX4uXIz6mcEiCly0gThZpxYDYqpHiy
I4hfVNHTOociFotoML7LvpkFPfTPNbaAt43d7sMxYF7wQ51nT6v0fsaQYjVmzOXLxHU6rLmvfBnp
iw8OiS9MfuDjh+/SoitBY2raAJfvJCp3FldE1k9k4F0s+2dkNIvOgn6FMfyRWqsJmc4eZbDDdJFP
IWWTJPNo5HXVoudvNoDiIkMrp+S2kxfswq4aC0ZTVkCLWHQOWHQ1z2id50Xb6TuxzIs2DII5uIAz
LUvmMkYzsOh3VUy+XGyZKBAJCP3witeLr232pYyMC77O9PxEqf7x03OOPYzFY0sllk21FRfLITbw
fgmqNIru/e7kyMzb7+l44S4UxybI6VPKxgGEQ8PFa/EIvU1/Ix6roVFNoiniIEEgAhBXeXXfan5H
rRjWDO2+jG84GWBjH9LGpmzBHj+GTuodO0C7Jtko6XzmhgsfMM/iAPCSdlg85ctW7xX6w3QaNZK9
qwFLCrLP5cpSrBZZWvHAe48VPxpLKh++t+6EpV9k7LSeHoUwRXe5u8opnmBNXpd57SL7Z5SC+8Xf
M+eOWQLJGSq6B3IAVZkMpnBJAVmIYjxIwHceAUTg6T7US3yMc8HAJn24xPbVOyBf7V8RbqlDyxrg
KQsv2I7UErQsHofecWTFMU2DYOnxcn/2R6bLQUmxkDrNAokVyLXPPMiQ/NGAaodNhfQ0ChREVUVk
j3zH+w7u9dH8l9XC832vuF/tkC3YF0mNVTHCUNJ9/4GdFJXrAJr6Np+ePTXeto5YLHproeMsaFzr
kzm4Y2jcqBuUMQTcEVaIBAoz413WQtAfjbNY1YbNBXgp3hFdPYZUW+fsmROSwsgsByXdR0/b3uc3
kTS7bG8EXMiHsGeQI5HcZKEsKdrSlYKTI4lKjApU9GbpAcOpTxAdGXJfMtgaM5x7fydb3jsM3M8b
nSkOew8BzSwcNx9fiR0NqiKh221EmL9vx314uFtXsPrAEo/LN/S2J8DbsWqUBitnTeh/JgImJXIo
/t4hE4qTGGxmj2/SGSuB7Ge3/ZiEFsD/hgxvAr6czhUDZxpj0f8BUxYSf8LEeqSXvwUah2CgxMPW
ZjMCBxXLt7Vbm9W2hFne5u5D9eWZvRahZitiE0S/rbhSFK3zL0ALSj6TqUePbzmSNiR2kGkeMcTW
WJWk1vyaTQkLktFkltFTmUHL2LrezDdKD0T9RIcu6d0x6KFMaabq5kxmSNDD7PnZxFRWgZ02+BJ3
XXFalWTb5AtjpjJslnuC/qjZxA9k4txDmMjmeCa2hSGNe1j6V3UerEDXE6VtRjsSEJKXXhcRXlpR
Rnf3p78gLZZQhKNxJ+6Y1D9iMlWjLbz+w8QUEzgq5UHs/udvMCTQf6MkxSOhzV5qBJdpQOYbsRZw
yYYi+DD8urPXZowzIxSgItoQ8mvRZB9jbAXVfe9C7LsKenfgfIPAUEQ6ehwkBmvHcur0wgZAibnl
SBH7WikOcfcpCIlvKuToX/hW7U4IjMfSzk1zBFSbGc5UBT5yIj7Nyd1UYP3UqjqmoJqUQ9HzRE9Y
S93ApUIYMG/z/by486thgWncJDCnFmWRrYex9ISqY3xij86dA4fYF5slAbnsa8MtR3HraQssZru+
aXIeOqcCO0H7zVS2B4fN7nqy47HNkqLXs1eXQ37eoHYjwWHw/oMoWHhuNGODGLyWwkK+SThbW98K
GGfl3ufV+b5Z90cznl0vNq7nMAY4Svl/ZvaNA91gzb1177ZEesm01XyIJpJ0kus1uSu9Khx0kbR1
ERPb7/1ODgHRHjf8HQRuVEGCx/YEcZ0oNTQgs+J+SMkd3yeQ+6PL/Jz60qfRAhsPFbMAApvB4OPc
Fs11xWaWEGzSUdz85g+/TZtnyo1AyDbSOOSdH2FYlprBi4lH5uBqK9wHeVbPDEIKKlgCP7/u2ilw
++vZwq+Iw7982tUvVrwEDSqbjDgzxVAyIG3C9B2lrvSjplao1mFFVeINPnqLbcmAWTyJFnkJtWaa
4kMug50wRrBJJ+jnAuNejWaALhk5YFUeFsxLL/VjvWexCFzanvI2SqmOwkC4leQsVNa7NOrXf8bO
1OhgA3VhD+1GTc5FSEqc85YBRCeFlw9XBxhXTy/j0oZe/qkKeJo+zt4aZAqCFuoTKRkV5ch7XPlf
esTkRzdX6SHLKaj3kfZ4ERCy00Z8CoXuS4re7eHmALCGlUIM4t2q5uil+lVsfJx6TOlMnMIb2K9w
LYjX0y3srrSjZC+paQf252GD46MMQkvV8WkBC1MsTbZcoq1emf6Lx6dNEW9RAd/ifUfGPHZPPdAK
zQO2JuHhwgBOFh8V5vL+KJXzs+aRkUlMvIR82nd2hfZU01YkZCOx13F4cGIbV+ED8lTyKMcufsXA
0t3Q5tjS/Zih8hrfvSAhe8CRy/BKx3SMtvGR2htarhLT7PV1JmYDUi/Vexn1PPRshoWDBpHjJmDn
4b0MgT6EQapVxEMbn8Wd7TGC42vOMJUVwF46oe+NTK3an2Pcot5Pkq7LX7gAOzTMrIBbnh3SVUvB
V1BLXzl49I7gDoX4gl3H78gJ9Y0/+OcPEQHPc6kuTnxDc1tZhfvm4ZhTNOeU3BipAECDhU6PrH6I
ScYPPFulgzlbjwIUhBAve5yDlfJE7EKrzxrZJDxdGHydQe6gdr/JC43m6TUe01tE0lI8Ae40aa78
SsvYjv0iR2PsRjcKuq4UeoqwnynvgVWNOd8Rged4XoOQv7dO1+BeAwNM1EgcLu3S5P+6kYHOFACD
cwkqETiB8aPQYk05koWoB88Mak8bkeyh0eq9Lx8SLOqAoiOx905/9Zl4C02B28kx37fFf0/rhbLB
gR9L8o15N3dgUcwnTerNjvRAlsuPIX3ntv4rWDOzY1+3NcwXRwvsug/iT8B58RF979VG4R3/ZK/N
va34FvUl3ttj9wOHtX0xfZKv4Z7BgX8KiXiTrDafeVWrnqJNJdRlrvwh96XDDeV9CJWGgHhT5PYF
4jnpcnfkd9zyOHMwJwaotqAizFeCreHGsbCf5ku0wRYCNlBl+kJbmkKLvqCSQCH6x+id28v4gizL
T8Wt5i9p51kvTrHhXk22xgcuKiEZDBnT78MnLsg/sQyc/OWjc06CksXY82nofaB2TTnjizBm4hiU
zUh4IgFu19dU0d0ZiERzPTZHePgE42bfeWOAdzW10dViOlIgT4GLr8tThIJIREWHsmQgGLotDh6v
GA8vScmrb83ZO59i4N/8g/NO6TVIZFnn0XNX64kRU1fB54vTdB558b5b84Z7irCMBRvTlt5Z5k2W
U/MwOhnWOWiYfPunwoC+xRSggpJa6qBXMM40wUERSw81fjutT35/VwdWdngzOigRPspWN1HOYX4k
SyZkPa6A0LOKi9Ux+QMQVmQsz/Xe2+3I1+4yJAiRwniu9FbFAn34RuMHhTdbPxoxIYC1kgO5fHFX
eI2i0EDgCMyb3hmxX824Fn8IVBnS5fxfm/ZtL9vnU3pXOmm7y6p6Vih/8FAlgq6oo3QprB6zMHcx
bcdB5gQtbQPJsLpBBnNUsDMKosKzz17JqoqjEdbINOCVOsJnwcJMZGHlWofFbRmU1nxJGgg1ASuF
kDaeZUJR4axL/0mEfBCBrAS+AhdppVWQDJPfwcD/DPjFbPrayoCQSegVAoN6O9KeqoDzTdf7JK3/
g+or56Ftpc84HmNo7iEZ6rBX5BOBDUwH/T4RF094TNA4gMOX+jCsS+Tt/nqzGkIWPxbpzpnEj4YH
GOaOOJFAuqIHWZBiophAHONktWLqf4uZbNhx3l4GVuVerZtP7TBu1s0lDBrg3KAijMVJsueLdWIV
YNi+qzOwUAoCTUG5/DKCn1dKTLgxguHg2Lu//sBSNcT6F/CHtOg3nm0JMsQfxnlBCC6nGV176qYM
sUz3b+BDvHS78xnrYvIfUuxXTKDWYwRDn7rYtaK6cwWXMyZNjG/cBedEME8/HyhjIxea9GX28tbO
OpJ30vzCTpOWz36WJjrtKUFzP9gmRqgWn/3MCtyoHvd3VXRB+Aw150DSbe1B5IEVXsmn+xT1uZqj
5ksyKEitZ+DzPWfWIGFvyQnIt/rt7Uhv6h1lBBXmO6b3R/ab+tK0kAUezwOew0aRRiVaomedfMOZ
U47nTN6CHN9gS46au3PJGQHhyBCfXaoyytrXDyKdYinGnBVQBY1rdrFIPcPnLadAtvYAXreXaICI
Zfn/jnhgFqvkggfKY58pxS56XUqxgjVviLQ61lo2WvvE5aUK/5oXDtzfuhgFzTQD0dr7D0huH7NL
K7phQj0HExPbktNl9C6tlrRs1CdlxaGRQSTjiCaL8pJ9LVMAMY0Sj8MC5A81iPagYfGyStHNQr4A
0QgYhOFSVE+27ULRKZCFO06cOXr0PVufG36WCkrCPtV7nLUUnRfdW4pfPqjKQiybU1SvcAoLveTC
WjLsR7ETpHybZ4PtG5+phHILUri9VsZUhaPharcuQ1E4VUTG0WaCDFMTn62uhosAfFWHslAtTNpX
tv2vBqjMWY+NtI9Pej0Lv5E553iZFz+ZCjikuTYqYm0PvyILyinkEiR0AFADCErvtRq9G8oVQrxO
oZk4ze0OK98zuEC4kd0y7nEOmyIWNbDRGWzOPzkRjqlij0/WGtG5206wJ2xvkguV0L1NEb6tms/i
lrJ5vdMpbDb63A1gajD7XcaHYC5nolqOMkzgVllgc1zCG5LukmCOUL/5hQ6UtyqzEzi0XvhZ4Nc3
QCqyPJECA2kMF050CxzLgH8+Uuc1pismEs99OAvAynXrjWuPTRGBuhLFc+/o5+rRM4lnG2KgHu7z
De7qSQhFdvSgcw/GlCWViBYKWIvulMByQdORq5mJanC3Habzey7biKbSGGV8AmaXw0LblWqfNoVD
w0joRdYZxXStPmFjHAwzakIyX9Kf1u3XCFoz8CPv/fMm0ynN0TfzZ9YdwV0iYkORkrTOm64R0viZ
pGr7DjP14VWib2CmfxzQLCMM/UwdhCz/s1jkbbPDbcBxw96+VDkVyzfciRiwp+tJ5y/johP5ZFm+
8rixzvTb7yXrl1KlYxUzvc142SWuG2jousGl8tV41AW9MliLDN+6MOGOBVw8LdzbgVh6GSBSye2N
Q54QhGb7lWY/bDaWwfxvzGFMTQU49U6IIYvZ4rJefCq0tImtXSLMsw5HQxadz/mNR2sX7s0Xwxh2
V1lvMYAEZUEA4aYyM7aEksmgu9NTxQF8mhKrFsMicd+FVBkPPaZTq9Vhha8hAqmmIdaC0mLzWbxQ
fP3iUvOLD2zlOQK1xXt3qkuW29QBFV2jQCaAK4gNVzuq28XGe1NP0k4Mc9n6EYFX0QYXo8MwGJwK
fPrsQCjLPG9mQE06KHa/aVZKLoVRbVDvtoCxouuhMjuVv8rMfm9skqivu1Kl4h5RqQ9NInW1W+0h
TJusT30eoMkYZ1+TFN2/2WH/pZdHlRHycnP4nh4watiZnC2prvETT5Fvl4kb+OrLtu3IiNrvr9Y1
BNo7OtBk4UIhT/UMUe1DK9wOr7RG9LpmIZGA0m3U2lMj1wuUp1sVC/IVTNzwOOruKH44WEVfgtus
AV0pR76prcyghdD6aepn/s9nv5PA02sXywjsu64+9lCLgiUehH3dbTRmIhjT0kFMrS6sP/wksfio
IYfGR7x6EETrrruAAEfAeejwzy6rbVWP22G0G+YmGqU6R60ZIZrM5OiDanHcan8rIn7S7gzXg5Y+
nCd9c5qrJcoqiXLIuyNs0SJq0ncfv4UPlMyQtCeO4z3P2TJndtmmqRaEHG3TQJoB59MQosvEQTPp
w3f55mmAK+tU+IlPIaxm8IYkRQ8Pp1yneg5p+0If6wMVTQ5zZ/XEejPYJz2VnMctgjDqutwZ05Xm
Q1MutqCO3tfARgQoSlmxSnnkaZmEBblXLSyRA06nUBAz1g3QUMMeEsppUR9i+7K2CgSzkSzAM6oE
U//oeaPEtDHsevX9iave1beRJ02u9tUkL4X/HfBDInSjZDovrXX/B8qXQ1rGycwu0GzbA4k6nung
8WRJ0W40T9bRNgDUiGGf8UdBQMWfcRVCxzvtioGTSsbxJAnnuZVVf+r2tMSaq2YEWMEJjIKh+tnl
2BBIxZ6EHC1ggSal8KmNhddAM4iH/yiCvDYhmFYBHnamANzzDEyMO8Li37YWwoOC/y41cDoFLraM
MSOcmmfz5OoYR6IYo+kjSOpDpYkrFp7HD32FEYdy5jVE5QJYm+0TwaDOxWrqrfqRQlIoDMD4UfKX
J27oYdv5dAV1Iinj47jGH2oT765+wcex/P0GqD+5850b1vxBUQwwAzWqxq6GqaOzmLkq9qW1Sn99
E9+1GcamijAp+Cn9t4r+TOPfV1ivEYRpNM5DoAR7XuUHnt57JmN/Ec16GHqIj5P/GG9YdiAl7NDl
DjGo7gPquJ9u+RysWACnu508oV8dznn0OG146j4ttbksth7T2aZOmTqEjZMXAikSKhr4MtniUcvT
OP7LAQQwP9fT8nUIJy8yooUFL6+hUK6a2mg+5NcYDiivPX5BiLUYygPeTeDC1XuneF4lfieZ3AQ/
XzDUwE8JU1GHJh6bO/9WVdiyilVamvHjXqzY2mDr6TRMvRts1XqdZ4LM10C5l/ybrI0B6pEB0r2b
38iFOK77/f1qFLQcuXurQH8N5mo4GfHeZStfoltDcA/J/TXhTql1Vh4fqKDveNy50GFuLQjPu5Mn
PGbvqiwlmdl6YuS0neOierF2VM7Ni2ruiexe4kZgb/bVjUpnO+5o5luMiCElzUpjlueW3Pup29RT
W6ofKRjZ5ozNayeGl+IJrhRJNpc9Z+0i0N08NMicvCGkxcE9crlnlNQiGFqCtkWj6yG9dijTvaVk
Uw46vhiC0zZE+X8Y62jBHYES/CuhflYa87tceoT/iKsBSBdoabqU84AR9FDf4TPIp7jlJLA1qcWb
mOjlVpYdKvLRKpbqa49B66Dbid0ZJkgGEePADz5ClXk3f3vApqrNnb6hdkiChCmpR94ziUacCvXz
dpBdf0poOPG3bP5dSaFE9NXwFJBJKoGLHsAabGFqFjaDMQ9Hnh8h5GibvBibxlB6NvScp4jsrtK3
2+Q4jzaQ5hMiLoyWg5KHDUR7bHsA985f9rJkIAqTbjefFgl37zc3l9654Fu30PcxEOkM7pZ/QQNR
CWAbS8tFUBKGwreb0Lwa/0V8fbrAnVd0mGVEC+05JmwJnxX9DDpTfxQT8NL4arOZRjdqy6CinF8p
vOS0NfowLbPejbbolJwQNV+iUT0GIn+kpkfm0wk7T/yMltnoiNmEsgfIryzbl/TptrXQMLbdAK1Y
6LqW6Vj0PMXRAlL+qbAvkmCfH5+ffVJmxK0TbI5BKrKwdYhOaa/sqVvhEW6OFMYQGL3XsQQ3gwb7
qww4K5y7uQ7FmDJ3HaszBbaKrk+hM0ToqrDDzUMcQclw7j1Mt/n3zpqbjVai9+r2KvNCbH2fwPMr
mHxRgtlpTU/W05+8CkclHbEE6yvpiaLxXZIif8c87wPr8Qtl4CgFouPvlD9FyBUYwzzNLy04k2X9
fR8qQFAHV7bpRf9ordh9JnYSR0ksEU5VW18IJ9krHKv1yCEdh1Bfdp+WZiTNqDdlFbkXvBrsc6iC
B+NUnM3uRRg/atghMHdDxvh85nPkwVxVIyFgN2+vH/Cks24nEwe+SorGOCxeoJh8ZiDeV6Fs1V8x
41xRPbf7AbTa/pb5TxRswKqT/WE9WodmN58RR2KUh1wHYwqYbYsn6dNF6FW5FzVrE6wztcNq8dsp
K5gs1TIsnwul4AoEduPCulfJd+sUg8dLDIetxGFRFE1SesofQT2xBkZEYwkugqLvXiXgZxXROY2d
yv2rokJkI8YHtpaDF42vSi4Mt68yQ/5dPOP6ROSMEwpR1egelvwA4qt5IHMAlzQyVR6/PAg+BOrl
aepiF4SZbEYYpdI/s8UkSI4O/JlXxRLV7+8okwPelf2mYAms8ZdbnDQ6j1PJ73+b3n/4q2VNKZh6
hbHk+E56rawTGlL63zmyhXkJiIeQ6R0xjZW81B3Qwq9L7oje1wiPKBvK1B7LBYYCsX56o3VOCSOC
PeTd5K9cpTnIvabkPqCdHhejoZh4hV8mr8Q/PHRL/HtFFnRj3Mo17ZIyn+6mMRkBx/WKnMetbor6
TFxFG8u8PtL1sfxQkL7GFQbMZikg5/S6CihkhA1d1IAjF3S0BBAt9FHxkMUEIQrNnre40isKNTHT
X3ZEgl+JBG4vAlgAUTkhdRCXNQvCkzv9nPG5n/FLITR3kZIHzHvuaI3CwYEo24U439stFVKTaADv
4UIYEF5gzlwHfdpFmAM/Df4Um17TOT8QYlJ36ixaN8GEuk4Z0Xpfpb6iOq/QTpd625LwmhJKBmBC
gneGd5UNGxyFDu7Hj6i2KhbvnL0A/QA/dDdqKjVo2AhnLibGd3EcKXi4/1kTO/Bwog9fUTXcdDJh
2wcRZNs99qFilNZ1nsfppoY5Tf+oNbMpKwVj8PT0fDNc+Jldmpo45nL9bG/TCTTUGDSUaUpzwsQo
apsG3oOHfJYoFy0hRfoDf5u87XQQ91QdFPnTP50JSU8AtKGt4U5U3BeT1EW2UYHwR2xfwMoqHGTU
wPfoXCRusLKfgmlA1w3xz/9p6yZ0Kx6CG3IKZgsEewlbAHTb2ztFU4L1susHpQYB/Qs5NLppiwT0
msrvv5JFLqrQKsA03EQzEJAgwoouLc0IPdm8AKLAu4ZRtguAn9u8Gl/tvKT0lpAAfSVrIXMNTwxq
rjmyKoQ6H+UB5KpTyysWLlCegIXMyYmZgUaDpCDVUR/csFJ9xhwM1Q67NE6icO3CzA3Grg3pVV61
IXec4akPE/oPIbiw7Juc9sGON3h+ollg4YUPoF4l0JFrL0NnxufeyCpBP9S4fdNwHoZ40sbKu3Qy
VctuFmuKshPvAKwVlbbdaoShEJ4503MCD6yVvAYLQkt6wZd66/ChpzI7XoXyt67qN+57daFdJnIX
DUJFndxHVjqaupYAua6uhO1yxhSZ5zgPt2/Y8X+Iek0ycqdbFhZCro9dDcJR7Cl0jRtX6mxLHsAB
PKDBiOxgNgNgIXKoiX8H6RFgNhMon0ZH+LBb0MYLC6HjU/uKk9v9euE+yA6EZpaM1q4ixP5jZIdc
r1XKFt4B0p8IxG8LdMsPGZpkGvv3+JenCV/tTJdatF00vsr1jQ7afRFSI7zzcWGVMuqXJBLNUw40
o1cbbvG/qAb2qFWTVRhT2HA8aWck9ew6hgWkcbe7NjzfmFZ6EXJfGl1q5HzZoIf2IcsqDP7cggI2
rLrUxJguyhVv9QU7CX4fXvz9PTuzAaz7bXzVO8Vuv5tUb6KbGu3msZEENncIH6ZXioLYRVS/UccF
po+mExP829KKeP8Xe6RlwDttz0HH4Yh8YnXvUvykCwt3FMQHS/568UKUJiPltxsRlu6M+6a0XEDj
T8xkxD0lPX1/ZAlrin29eTKaA+Q8rhjGROMCNC5zGCiKY+sKHlP26btmMoOcoPa1I5ESvbsU3ToH
zhe7M5ZFELYkfyEoHNEQFWgdLTQcDnF105HX65P86oXCx90I2uLzhVv62IYdXiUqmESy4/euWlHk
Y2c/RxdS7jn/1l5NjiukynAOC4mAvCgiXfzNrY0gd6x2Zme3XfKVpxja6gITZLfJS1SmdsqHRF+l
G9Ut+Otk0jmXAPasyhLV+tNh2WtMaLkzlQQY2X8961iynYOAIo7RXeFuN9VBZVFLHLyxc4hLez5P
yhuSZlWclc7y++iN0/oxSCImQB/POeabs/yKNXnKKdDrAx7HN7VepUwcsriJ5P8mjoNaTas6R1Yn
0AFtvdyNUBVjZaurzek7CGUnG+kR8KsX2iLxd34BMHXmgTeKv//v4+Xrdry+Rl2KghfohbzP4+US
t6yQhlSM1eUJnl9a+9dqis4jaBMkhdMxof2P4xpt8bfEuiZy3+nruLCnWXTBXYJXoKDsUaprAFSy
N3vQXvvacIA1Vy1TUlcQPTNI/D5vnS5hqlsBSAAKMoj76xvg8hxI3yU2AaKOE5hjn8h/QexOu7cn
Mz71QrRBq66yRaipl/3rkQ4/CiBZvWbF+IeuAkilJR84KLaHCmsfgHLtkrwL9odYnuxgdUfGDXDl
SAZ49jK6svxhLPW0piK6zUCJrFDVD1qA+BxnRPt0yFx3ASImMlqqQOGRhcxtnAiAUBVAiJOE4kyj
u5+NkG/CyhmWIjouSIWOEEVn9xlS9DpnF1Bqzi2p2siiQNsM8QqlvuzhY8tobpO+wHa11xK/QHlE
PWD8Q0XteW3l+FYiJ9Pwh+hEGJbzD2m6o2YGDQRpOMS/99apxefGtGI4+7S1n68XkUJNcQ+3rNB6
gG2XRQ7l1MVlSGH2Q8UPnIAj7TzSawFPob//JN2U3htt0En/IQJIk2KDTlZjl3Peq4O9ivLGj92j
wczZ+BnjhRA8CPwqqJwSqIwc0dk6HnboDKIwswYuUksSJjebUuS+BY7LvWRE9rtj6edHzcac94Lh
3rjInXfUs+Uw6pcZy4fO+rM4e2I6yG7g8KHNraO5ePvExeHKoSMRGs1S4/5syN9iHFp+ogJYIyrC
2zwuG4Jb26us2rUJ2zqn11gXegUSFAONcavB4O1UPzxjkqHVl3hzfqAjUZq64OmvVwRJmTnbHZr/
6b89QOcWJEnIh7IiuiCkN2PXgSwrt35v57wHalOcWBYLbk5WdWwyvyi92mNYrBhtKWZ7wD8bjPoz
+AHO/FZ8xpRrf4xmZLhVPXPPMc1Izj+foTkKEmkEpEIOygGQL9Qqiv3wrtsCw/QIM6/KBBL5Twrn
4B6sOVwXW8fe1r80Pwr99vGxPz9IyztAsTU4+J/7yo+3zeU0ySG5FPZdCEprjxGmFjuwXdEIdOk8
yfLN8SiWIz6UVWVQuvfg6jGkKPrWgW/+qRJ9botH+DWQcwRZ3Z7qEel8k/lkqXAikmZBOkA03V5T
wQw9iz+3JgCNAV9qtES7oIRBFvwCLTlAUp5o7d2sUT1JlvrvYbRK5Myl3voN5oPkuh+LGi4sUhcQ
G7jvq0NHP7NJ/olB7vsaPrYD+lWMWsJsn5jywFEbFy2+RCI8ogcTcXwsbt31V8iWzpi+Gh/sYQvP
jfCSJDKNdh7xQL/ZgoRMSQ3F71vbAikDRzQp4tzRfQcYSOosgPfh+EpGR+p4K83Qej1elRyQygAY
IDzZ+buVhkpFVslHlsyuP7MvLRqBC95Uycaai6DvL0tGu6vjMSMO01EKOvKXyVWj96MvYZgPL2Aj
cqj6teim953Ioqo7GJe55wECRFfrw53eIe9ZVqFKCZ65s+E+VRLrAfoEnJqNQ5PPjForY8AMBHu0
kcatiuSdd5EQXH9BRQRK3Tpisussm5dZYg9XKklL8gXSqJuZH187FAwVQbIGDeJfwriTcHyFHpmQ
zpRCjP7l0vPqUWGNUWeEBjuAtr2PGOgnohnQ0Ed5pg2uz8Vyp7OiIEtw+ZortMjuoGDohlOIpU0s
Z0S0pfBlkUgm2Vq++1wXRBHM0W9hCbhzJwjJ92QWYl6N31FAiiQ+Sq4iGF+T9DSKd1LEBOLnukWI
T05wGwiy+X8ViZtTavNozcuTtdHbsrrcuA2DSwoi+AuPoMAmutxR76U6BdAmpPlyxgLLsND02hEf
69EJYSC55PpIAuNmhbzCKD6njBhb0VbqaVOsvc4KntBDHrFuhGHoAxrhcXaIZLW+5JouYcPmfmYs
EPjTfKc0hlAdgdZyCFtWGu76F5M47V42PHVn/RVEbO1poSffSJgupzhmrdrOGNpRCIwkzABer4hT
1pwpd/hVXBt3x1+8JEhA8oQ7IhZtreb0n7jtACbiG93sUDJlLJp85nJwyhNC2r5JuPXmBg6Sa8SR
Y4zirHHC9R0WpTiR7UBa/Sj77ve5bsvANA0nxE20cSJhUJYNHdZKQhVGINr0knBDfNZNIFzAoENG
I/Ki/oa6g0mpFof73uQ2Z0WBiGTYTpfTm9o+MHB3amn7GqNtRn2qrC9P76yp7yHjmnm7CreP0q1a
+S8gtQhJh1ObISl3xwm/GnwA2tsuZ8sofHmF6qR+ZR3hwr3mfeM5fjXsxrXZb9sA9kp8dnY3NimV
g7+n9mwvH1Sfpl0OLTZy7IR1CgAruaCxGldYdxCE5xbcvFwpWU7LcYv/QKialnhhRuWrPi92wBR4
fO4LYa7joEWuT7d2IqMn7VaHEGay7NCd77ZZZhj8BOKtxsPTHfeOrVshLKxfElcdk3vAXWC/cYzg
RNoJT04Vu8hu2MiAkN+zgACQygSn5HKofJG7GKT5PikKy/waf+wGOW2ZALjBP1WdH1l1Sjj2yvSj
slXYlzsr3FzEnTULVtJ3LjMPVQfSsZDsL8yS3ax2+j9r9NrTPZ1WZTyQgzqzpBsCLVsOmtEjzXB8
3QXDtssfxUtAEuTfs7ddjalal9fj6dqcbsFnxyF0kFF9v6ut0LaapTxAM2lqqo0JM8LpPMDtU4WK
O2gONFU1xDsjTqCUyp3SPr95Ll4iqYBzvFnIKLl2XBt2RpoyeH49yPQDdjZx03HVpi9vJF4wAfM8
F+VXYZcZQd3yi2kqMC/pJ3CeFLWu+9j8Fq4AgY7uduqOj3QQaiVWM+h+AUFomj+g3Qv8jUTidRBW
NVASmFEXBr+MV+bVs5oux6h3bqHxgJoOLWxn0jZH9kDZ67RuyyufAJ0n0hl9c0FmVtL4BG0TFACa
aXafrhxiclwOqSrg+SqOblE6qeM3wj2f3RFby/WAU81iTeTEh6X7naywGPaRXqtYhe38asnYWFYG
X1jNeOzTptokquNB7IX1U+AVrgN1ld4g2hX1I+x9Umf08sPdGrEFBbMZfXZI0u5ktICXDeyW3Qv0
7jF7kWOoXbo7Nhpqk9Zso4Y01c1xx8TqnffnScPUIyRzKOv5hu0okLS5+ilEIZhgUcRTPmSO3MIh
9VvBnwxTQJ4ORWHGL5/0HRuWje9DvGOD8XWVBzYKwPY8Tx8M++tfvGXVI7nRLnpB5dQFqetrwb6K
LATDVoEG+JMf27qwG7W0eyr5WM8B28GptoGMxOMXDwFgyfIMSXOjSYkykPeAwCV3tK64cziQMQl6
dpSViLC/Phj8KoS64u7wDf46JuzIEvJ36YpZ9NI8VHOKIRuCUI5dKKy1NIFOkE7bf2VQDvGDPz66
NvWWLUca/2zuLtzyHss5OonXQtwN5oqXD4Xp7p56vuzklQY93z0ntbAHOyMFxjByinU/N3zhqrkG
bHg5qNIahVcPDMx0yo4/JfoKD7vo2s13Vq6HM0+a349R2x1ourwLyew09MdmxcrLpIn1dIT87q80
91V1yZ3IRei3AD1NJDt/QIGeJsuPtz8t4UVm3jlqNH0Dg9imgQh2xgkxOcjBpPL/PJEZmMbmkS/R
UOtJLr4yr50wv07gLeDP99rJTb7hMbVCsaiKrZEv3yt/AWEo6LV1kD0pE+49Qf8UBUnWgV4bUVzq
6t4RtlpVAIk7hrRQObs7EuwszA0YFRPzB31KHvskUo0/ktiY4J5DQfvWxsAl1fI1HAmEmRLz2tnv
ypN6wHj/dbvsO2oLfRDBKRSjqCqjnma4UMg8nsXO7f2ERC40CWUCNZ+6W2U88g3GSgHIlntRI9Ng
RpyLXsBHqjmOnTwZCRvxmyJyQ5rPATE7qZE3/P6+NnljgOt5WI4uSHkgqpgSfKyu4WFpdcJpZsek
zLvQdcZLyrk9MaRmwRH51nr7DPW32ZujdpPKTw5+R2tPpObgQRA2ZCsWKJ9vXVfwzBnxZhLyLh6w
RrTOGYqhxroLPHQSXHPNC6FpSJMA3YvF/jh8kdnaWk3N3cebrU6LmOCfPJ3/qxHVHyhjJ8eH7Is9
HWh0Ye2ThsFNskgUphOvQsq4se/bxsL4oemNF0hSSVzM6cv0Ou8aAC4x9a1ULBqdDJ68Btwh1UCx
+fAIDY1OEqAKyOVY8D9A+rnvi204RjvUj64eb5iZDU+UqVM6VTAH0P3D4tq2lLSSLuiH83koQox+
RWg2JHT70/iT5Ux4fjwHrXnOMpjPdHb3h2QOQOUAHEfImADV6oBr/OIpeyJlt8R+7y1NlscXXbiU
ZOtmgJis0wtWIdcYI2EBskSk8AvAs6m+MZ1QhguPdNyRcAGaK5GOk1R66H+Ea01UG0E8btpXg6T2
pGHlrk+QA1/rPkE2VFsUG+9s1Dtmu0DJisZCCx5IK7tZfWZ9Nb5ThZ7xa3bTR++S0YRBkVMomIRz
KqWrjT3He0ac8zzf1VWQbGofC1YlG6dnW1eGdRW5Ha6SKcGNpOqoNWhIsjkkLPkWRgzQc0rs5f5r
oUVmBS5ihO41BYxUQmgNAcJz+XTjhjTlLOpgLyjsJIf23/6REYgzYhC0cG5Uk3UaOyyONtD4i8sa
U8VNpmaw5ioDhtXh0webQJq95yS/2Ekvv9NCIJkeA/cfGTUcu5koHmX4EAu50mCMB9xPJDrXji1h
+8bsh0tQa2zg68AlP5Sho6kCERGGSL1sAYCPWY+/fZeCenXAGP0NgxGtXVP1vfl5AGTnEFkZyX/U
GbCtVJbTaLVZRxQFl8Q0m0Hxww09PyboLaOZqYnnC9jq55VyKWT8VzE0AiVHShLMPIsSRCP78UjQ
zlRdnc304QE7Q2PYEyaYTac3d96DQ8nQuXkNYndQSKIhqttGgLGG+WtFKNNp1kHpB+GZdeIae3HG
Pq27/WZS7CHcp5mK7dUV+qXBeiNuybLSm5XzoGOd4m9HcymTn9VOtr0fo6fa9snF7mrASJbU5OAx
EjF4t4XIBl7rcrWyojV6GXIdDc+64F7U0+R1y4DTnxIkIVztazIt90xtHI8PGb/uiCjUqqNYm/Lz
PsXFHYmuRIcIapNrlozgmgLnwZu0Pl9iz+/qIFbSdAUQ1Czfd2DYunUjKS5ck4M1WuasEi0BPaXz
+/XjMBWiqNpUS+dZ/88Nj7SzOMsCb0rBKLK5NiFDrucSzY0NUVdepn8aLQB+2w26tzdBS48ObfWh
zSqfYrGgN2v8ydTrIG70b+EKt/7ybPfdP/8FJx9SPN/Ar11i6yGjmwgktDg6D/6tac2OW8O6jh43
ZVT27WifplmyIDx1iKD6LZOwpWTT2t99rswEWnB75Wr+3z+Y/4T/tthPrlZaLInO0wVExAtRu2N0
sOuQbOj0Hv4SigVjyOWXQPkVlJw/lg06SVqjpYcrHrsDTMtarGkN8fBZX1yUf1GCLRe4wfhFrWAY
w/KpZkHLuG+rWzLmEwwDKnuNJ37yqnwWlQzCAse4QE3i0ZSyQgyvs3rm/uO6anBOpJiegXveWTXQ
aOtai/ieaV6U4oOriZeTRkVuXofm7d0cEKs3GHQXM4zjrXBv+A8JvEYVYi1XzmyqurLzMDY97vkK
Hz841peHnCCp2vfu6N3d8EXaU+pc+LQLGim1pVdMgwak5ghuKfDx+XrZPvvpb+xxm/fBE0Vke4qo
eP2l1A5x31NYFRqgnNbew1zXx+4Qi59Mie3TB29YrPa8CK2vvJKO+P2T1SfrleJVV0kgTgW460wX
upAJvDQJ0BIfdYzUF3eXSUPxaXmMszpteumGqoEnvQcg+WVe8pIDY9Yd+yuPh7Wto/c2U9dcbryT
pcJ6JXdMnjW4XktiYqEJE9/u+uat3ZWrZNH79a9tRh9/j6dN3htJav3D8TdGx7+4Lead+Gzrty4z
WUM5LGPBZvIFaW+YiUhF1V8aKIgQxW64tRmWOeYD0iIFguftp3vsiLpyz+I0lyg4WEdssnXHpGT+
0jV3U4iM2flXZjaWzD3LacQbkJCGbm2G5rHlLemOoBS8BgzLOL1qwlVEP7Hh0jOYsdW4WJwd7ZrZ
yJsJcIaPD4ht8Y3fB0vrmNStQiL34RAhE+/4a7i0HvS1TAnPe4mfoWrEf9SlQGbEq2UfGEXxWPDE
vrZ5bIDnIMByQ/VTiomnSK3PlGc6MLKKaKeY/UxyU8gRrcdCZ1RIiuC8mmRKKKTjkrMHbwju2wWZ
jQ7cI2Rqe4oYwfl/Jv+vXjFGJRma+bKmbaV4f4LVFYNobb46pMM77V77zmaWo7m4flXAp2LKX5nk
6LK8Lk62rQ6EmAYUbkXh6b8//uiayE6OJkF1Ze1z+us5c+yMlOYkEdwidCJ1abBUbRtCKI6TcPKY
K1JGpTOUJeTHu+tXsbe3xGKfiCriR7Fbm2/354vK4Ur7/4YR6gj3vJJjlh5P7KESK3mhm9hcmBxh
3Z9npJHf3Iw0t+QzjhvrmSZgp93/vDYutFdi8dTOzCbwaxV+ozhKuU9KD8ht0jfeaZGDpmix7R+R
+8eX4Mfa7DExlYAQbTIC1yX6RBe2sMaxNgkem8JBEaLfpZghF/k5fhY/+nhQ3rtfHs10zYqmjwqA
rsET/5wNSgWMbTAmW9XA6mwlP0kOHakDLl8jx1bmSHROEwXje4L4PLJsYdGpgBGkJgUwfoRKjZ8m
3O0tsxw+CnHHUhOoxjK9E3WV3EqQoJ6JlbpmyuDMUyIhThO4HuyblRSQ5XYNVvNlCyA2qOq8zkHN
Vm9gSy7Ad7dK4q3ijEohSGYaIxRn1UcO5iZZx0cIOepKPKdWwW++i+d8XxiFFgGbyofTdi3ikRIN
SBelxLCvMOf1whusOdZvMbbtzg18LxyLrIsRvwT2ScnhZAMfXdDXFa33tuqA2aAbPpUGeRh6aKQd
9qSklf/NdyUY5B2D8frjHxcD8/yrQtS6n2mq71+yawoNka+8xCgIKTtQ5AJFcF7LqTvrpkUwDxrG
fxSiDbEIxa4ANgcd/WC06rMi34uparVUNi7vvszNJniki7WUee03mfoAIExgsyUKCc46vMXUGIFY
bzO6pq3HzkELKuQev41lbS8a77vUGPH9wj+ET8jlY2QqHbKieucebLyU0ADrdmIHk5o1FpISABZO
38hht/xpjQ0SowuvPYfvnJL8ArFmw/Qgk/8/d2Gz5oOr6PWsCez/lPFH/LQkMgmYWfz95Sftikwm
BG8hIljamM2E2A4XjlIiGOigT9gJ8yhXcOGQwj8r+3jkgXsCQcU8ApH+KinVkSqcx+I2efSAu+ul
8DhGnV6XIWf0pI84UVnZ3lGwhjkMt4TrLUbN+2kjnBff8wGU3OQ5yzJ2b6PGDQ9a6FnH84oFTdR6
NWaCh4q/d7gRICeAVEtu2u93Yl3fwVDtBd3C4FFlIKM26aGgdijBluHGejP1azcCVJE/3q9z2OlZ
Fo117LKN7LAFGx083GXFaNKM3qfjjYLtvxX0hlaoKX+1/ZwkcPxsaVVMXBp3IioTE2vgX7KTFySl
e2wUZX43/8MFxS8yADLly4BH3J9NXKfFZpRupnazxbiV/JD7560FPReWNkpkzZ7z978YAcM+5ZFD
yrXBl1pdMxLSdMrJuvZ0mmsP43uynv7aW8183nZWYGP0tyZPsD3cnEk513ttYPqRzzaMXyj+hudw
gh+xVQJ4UvmshFdt1Z0J7/U8bRQg62QWq+Zg2MGpoVWh4shk355bCrVvktdOfS2LViOFcrNAm4+N
Rc0EzjhbqrrUgnl2ILeczJvHpTcE1v0wWUTlcadgSM8JXhfczQfgXPGx5djZnNb5cqAM+IJY+Ye2
/T+ImN9flceJzO0sG888rRehpPgrJWjPQTkxP7OEFvcQKW1Zf7k6Sly47Jz9cMdVEy+xbEVgtMHI
9vN/gRbGTPtDNR3Zb+0uVk56atUrsXPqp7l/n5MQwaaraaKe565UXkpWMTHsYnB1z+bam3qGPNAW
TuNiTAt7DVg3lWTJFZqNwGVQdy1UHUzJtp/zzMRoCyYHDT11NmjidbupmjR23NiJerLoKwVWfZ44
jUw6a6SSpuomyUO0nt7M8j997CmEMjWInP40BIwcmZNtNbOCsqVlHxPsdxk0IXKFUe55pR0WAHjC
Hl1q2uEWt4NoQFXa7tjNAlcCVwt/Yaf1PSZmNO7ilPDW7UDSNAD62CPcAlIK1xNx8pj7+BH6Q/vt
4DpZg6s6/qITGCj9Nuy51CoTik5p04ThFbYIZK1wHnxkZzehN3yMpuE+8ZuunJo8RCJPYTetqIi0
z837iglYLHhxt5jqBrnseGoEyeWqNpx3Uzw7JnKnBqJWgn9s2chUarenVjNxaS1l/g1BW8AcvHsG
FIlqjXD6IZT5u4tw355BqE60HhVpMIozUw9fH0/EkY2RSZbDoZeXWMCYOHAsAPYYUtKmCZ0JKmjz
fIBhEPz+FJoYC0aYSfgiRcW2cxNCAeNRpCXrF8+XeucPKwK8fZfhDQrNaS5jIlH4m3apxEE2zsN6
QiLgy2VbOG5hrb4NsTc/EiTVc9nwFLdW+BZY6TaGmqF1GfVcnUlWe8FhSUy9zGgrocMnBcp5NMsP
+/x7JAT2FVHT93pzR3ciTjB2XM2WEObqK0t/z1LrRycIunvkxURteL/+WIdJB3uxSTuvhQJVE8bm
cQpo5UB1ttxkhY3qU9YWL29XYjsQMGDKnY7kn+UkRpG2xKdYK4J82TzWR+tD1k57E1Pidn0QiXfc
BxXouWzjVfGwtkSqLiSIWlkY5UdLBW84//GiwMlfWyEAkWWABeg/MCJTmxBZkFnPcQyy/EQB3vcC
d0tnHrVxtA2Ijmx4tayBIsBMa+/576/3QvzwLpoE1sdktVUZ29NM2a6+DrMi8oaf6aWy0BFasj6W
n8Rtxi3ZdDR0KFU4iLVQzRrNHPBv1saSyXhWyZ5NWmasTmaO3E46RPk0jd1WMn/AjlrTKEg1hNk9
RtJxzkPLcrW+QF71TVW+O0CSWo8o43d7C3rz6l3NMEoQzGoXfdE9U4N/hglANa5XURy6/GsySa7x
k89G/3FDsN80x6iM02MHkf+/TSL7c/UdzJe+Ky/jcByHs970Bq2tJX2QzSbqxqG2hVhRvPvEuV9+
CrmaNZPGEv+YjnhLui07vC9w/VdWRtzjpubDu63yctRlqaLiDiW8z5C6YeOUq5S3sOQh+j5nIATv
FCvHSDyUaeNerFdZ1WwdGvD4CeB987hKiMr9kweVditCQgZSP+xmV9r/DUjtH20N8BswKZ4heLDU
HoCM+wCDYY6xBBsWZAF8/zGNCRGGgrpUz75L34nASJ7h4HNW9hdpHSuHwxJIMAWs1xiD0mYSFEJA
dgygdHA++ZoAXIA+JAMzlqWgvHQjdoKv6Hxo5HSExyBEjoYhVqSKvMOg43uUNLNcyEVXf3Ee3cqC
3oG4RXC7/YSc01tcRKzarFqg3We19AJsFfNbT54ZE8BhdS7Gj9lIqYWgrCshx8jHmkQWIJgMFC9i
PfEDZOrrvXrVNbcQYCAc4Cnaz8n3/Olj3ONkK6JX6lQoMnDRSKN2UeRbUCeHgP45YWShBdz2oA93
bXJ4FFyWJwzwwpDuQzg9e/l+NhIoUmQwLLQ2bury1sVj/ctIwD+LMZRZsdV1w2cUvR6X0QK/f9Y6
/1LPXVjBnuyiL7lzIU9ieREMMltYTAQhBEbEllFjPY4rpcvQbasZ8QbEzU1F/64KdBq08fuBvVOT
Z+gq+BlJNNvV6Lo1TE7pdBHnhrTY7d/LqM4r+JR9YSSMayQHXQMEPfeRNQyjZBg6SrSUavFktvf8
ddWzwhLqJvarZwD23Bvi/G1d+WpIHdJ8IxSwCz6II3g/HBdiWcW5Pju0jLeVStGfbrCgnAKD3vyH
D0nZhY5JbtKWIs0oX5bKY8eejrMXOJLeZsAzg3I7P0IsnDD0qwXw+JJeoIrKz0Vf5x7NxB2EysRI
EVeG5qyfoXa/l5pXIA71L5s9SFkymjd8jwLjbZKPBkPp+vWrKQ2bNpdy1hOFRPRnJtWmug2FIXna
N1H38Cr4EwNMwnBzpeqWCVPRzhOCdnb5Ce0HVsIbRZmyX4cmY044BNUP7FfCjsTbDySXdmVpCcIs
fPrpdnzaaWFCaWgD5H1+0POSdxUeV/RsbK/gxQJQZ5VTHMoSO4xA5g7iKwUun4hMI8zEFWYFf1cW
BHyPvziJLI2zWL7eKN+C6r0NQiyyyQykUFKASBWdwk0Eub5W2h+79dXOPyQOKZ5kLIUbJEcWWXJo
OFIPiuPzTGmN88rMPETLvaki22I3citxSvUWYKTXpw0/PDRlV9nm4Ok0xrETj91Td2TKgPd1ZG/f
2k2IOJMg0ofsKBJ+mzR1SsXcl3VUWGq5hDWT3GQNseBTeKP41bqB6GTB3UBJ0RdqOpYYTnbcpsKO
e6fM5Zq9StwQeLQ0MQsgnZ7P5oz/OBHoReCsDoQQ5b/IFNmNDYjT8TXFCYjR95RMT5i2PRM09RoA
SU8gs2bcn/Q+iEen1ZpuCM+zg2/BQqGzALCL5mOs5sWdtIHnlbbYZWyQmo5bPhfclqqZPQ0sUCk2
YJeHOliPj/vojRJpZlW66HaSRsxibGfcqQos9ewcHBacvr5MKlAnRHNtaHjtuVQnani/WzwDwHqw
EP4rnLmyy13ZayflHVRsT0isQs5SPRSG/BW2d7r2BOD8SkT8Jgm2LzeK1d0a8hGUC4XzTkmjw/50
42HGrDUuzzbUxIzWFJKAIlvEjOj6uDDahOjpFk8xpPkBMXanjVPk5CflaOQIxqUeoUA4BSvqDZ05
EzXHBzeuk1LuLJx5h0bmG42mLJ4H0MyFb7zormv5Yvh7xArbh5b6bs1tDwTruPhv3CMOPwajXjhL
2OlVNg6kAaXMInPyPqmgbpOPh8Th9L4RSh3BdqCgAcKIPzACkrA9/J8RvedmhOwl8D+uqpjvW8s6
L46GAe+lxNoMRrU/AMY/dAN9pH9x3CYii4B4SEuFmRDLjJIaCogR7JmZtsUjTPfkK9O1RuS+doof
2rmT/maKoUatQg2icAB0Ev3kEDg08LVAjvC2ZdtlXy2S5T0hHtu2YYmKoK97gm5OQ2L/FhSAI3yR
6swvZy0SCH76s/Ih/6U742Phr5/zPVXO3cZnTyRiOG3SqGL6PPq/RVv4uRy2wlOZx1UjZh3Dzik3
Ks/E06C1p6SM1al6PZoiERTBsHcHIwUKNDoxJcdR5bY+FcgaxEdD2dc91138g+lXSMLrFvYZslU9
aoHbifyc5MYtTboJ5b88vDnOBCY5KnfwemMUoEdhSJJeRF7Dumn5drqp0JdG1mNihhMQs4MppL5p
YgkCAXutQW/ducBC7i47dyaQApRCWUku+ppFuYI5SoZ7bmZF2E/SBa2kXPuzhClFQqCkF/R0SYzF
vSC+TLY6273B+MIh4X0gxu0zmADlOogWaEW+NHYfYkC2lfXQVt9N6nrfxadSWEfyWr9qfDvHJi1r
uNaCU1kPY/R2l94sGjLiru+fa52y+6fIRhHu6hNBUFdf+6Z7JpURhHodeVT5imnY3/WAyAbTRGiB
WJEttLHGOzVJ2WOAun95z/UgHCQIYdlPhiMfuR5VFlA2ENxameP+6X2aSz2OPITBiQjVOjNzKSBc
EvEBdwPjs29FWReqJPmzM5xthRDAHGgUv4v5v7eYmgF10hNIJni5bz1yMrxyUF1ZJDC2FSV1019y
YXgTBMATeqsYDSZPndu2RrnS4AF01B+sri6y2Ez3cwVZKOmufZHaPCugBLgVvtJlcN32w5zJQ4DU
/bW/YuKgPcrSdTQ+1ruudtkfn02HtXpI3Izt6Kbqw3e954JKOPkNYlMzI+N0u7bbnijMmDsCZpbb
g+bCzMMHFlIGpWNWb/S6VQ1IxCn71GDVcNNcww0ytHmgUpgdx96WqesEz5ewm8cMq1n8EU7+utaq
5ek1h0qwXkDMvCEH76cyjExt3YIbQ3n4tuMDbLodI6cGBokOG3r6ZLcgQWTIGhXXhpiTw4NNbZYi
VBetCP4pM81RhcNA+hrnce+limlPrAqAzYreEkWSQ4kgVBc7qOtjNiulaaoWTBkRLRtGwN7U5OLW
RKEpEfE2OE+a7yEfacMBMcHT7gdY898nL3OsrNx72ATkq/PFUn//ooTRWp8XkDweMOrTCT7WuaO2
Oo3vP5rsxsOxu26cZ6Nb8Ko+/fr+VRczwESzhvMXyzsA3WM1jqbmCEzklhTJK7lUoGkI7iniSanl
UMLeRm0NVspFo/zUwAT53lz9vnsKI8CiOjCRTRjhJAyouMt70s/ED91Y0CsXWAzNNss02Yl9Aboj
lfWx1EtHYQa7zGz1pgIDXcBoaiYlvqsG7hiUfKW3lkalngpo6E76nDeLRRm+UwjUtpzSIpq9PBmX
kiTQ6B9NVssS5jI04G6QGPuAxNH2pIlX+ZVJq66aj5Je4WFOMt1mfZnIKYY7b3LxRj9YC0nHW6iP
cUoFZfJ0NVnaet1glpRR8bugkaML3ap98Xc4I1djmMGHAaVdlSvboVdmTU7RTus0nN4r3QsTaSWe
XOaB+q11DltIUD8N7i8W1gPFXL5I/P8SJ1Bzxr3u6k5bUYkwPgubnnyMoCnqh2HDTonETMY0EzMd
MyIhFcfjt4m/XNffzfVrlUBVR5YWGcYrhnVjy/BYbaWV8ceqAKhRXZcQ2oGrLe3i87TOo63EbsdR
EdxMnWTAxo+XfwWLKFGGQpY81SmNl7Byb7JlFOxMwg9MCT7dphTwrlh8D0BlglCVhw7li8Ndj/r7
QewlLKMSTDzMLkZv72/Ma8Lkg2LY9m5GNf0qU4cu8HZC6Wqht9g/zEz/8kuH6JlmgPy4O69f5DUW
KdVfzEJGb3tUne6fl/YWvQEs3i53NgnvcvKktmUJUWBYX7NHGGYmVriCk4ThEwhDu2vgY57b7oev
uqzR/9zloBmt7TsL6e2sKLzOeYbsDortvureWmGmfF1Op8iW7WdeY6m+hdkVAQ4qZsjyUkKLkopn
ePnWxJ6c+MnFwRSHWIjiS43CsbhYkrUl33v6MA36/sx1Gd/iJ7cb3by+u0cbS7BAC1KSDZwravrO
B0yznZpLScheJS6qCpKmikegYwj067Rjfd9OBywNfZnWSKOqUWeJrGPW5tbX2GujNf9s3joBqh1v
cgWS8KSa2xB19sokQRfQ55icpVRMKnlqIRyDm6HHgg7KVenrDeHnndMlx6mzKi5iM/7r4maeEbUa
LGO9kQS41nv+0eiOMoxZM48HWD4UvWmrTP3T7qfkjb4T/sRwtV59S3bL6yR9fqgVXT3zWlbveCDC
ccYEtVHHjR+0ugFBGpBVSRDf3ufP43ZNs2Rg9XkvI2zn72PCh0Sb++4Bs8D8SUpP2Dw/FHdpsaVi
IwhfTG/ZGAYFWe2fL35bEcL7wYVpg2cD7iQU6nUNcpWx1f92XsdmWOYOvaapKBQeycpwztk1IgME
ZqbrkeFjfrvwpJgHMxnLsDZmUW7aeG37leMhYAFxKh8lp+RGVR2zavakpO3dRVxDbjdsniCr3KZM
Mf1E3z4aPXuQ+oQgabIe9noM3hz/pfvVPPMwU/o84O2Ve/RL+/i9AVWaxI1+w6ag/ldzqaDRDxQN
XZkxtueZAvKrgUSwXd0ty0Cm1eJQ40sgjzysgEvPvV5imNYnuWEhjBFdp6cr3DU1LJRNLaBYg82q
WAa+1ilyN6yoHMirVt/0nwfdCD0QaLtrFEq8yxsB+9KDt2LURZWltcbrf47dDym64BLNGpMNalXO
SokKTpZhRYUejk8hEccY2Yga2ak1VfSIb2ILCp9G2JcHWCw0bOryW7k+GGWwVbPob0V89O3T25xX
fEAml0UC31HfMNIjIGEOOsdWs7FNd0vdRAN4K5mmRA4IbnjHQFIyilR3gfJetRzJCN+oZtbhTJD9
PGswf7qkMN0fTCQcJwWw+ifIk5IDHokCNZzKpZatT7rwBb+RvDIJk1qrZjSRGwEKdH7EsdevScGU
miUgk8QQ6nP1RMHPC/zPKHzG+Z1zlNeqWs9JQXQXYTJdgNF4BW32Twc31x0oJxNiPXZPTPzBUBS5
OVQQ+2+scrGHut55+mDMiUjnYdZ1f5wCyes1i8WM/lMDhUncVDw4lPYnLeDPTetpfUFocR51bOPV
f63phIe6buCbDDgOMgg2DeUoh3qfxw5jMeekdA0Eokhrn0prPVSTm0YayzIOEk3VMdRB4Vnw0Cz/
KbDAZhgXaeoZfMIeG7WnIsFI5sAy6FTpBVfCcN8de6JOSB0xmaI9XsPoE1gCa/Ilz5dw/Ftpty1r
BJw24rwd47j6UeYwYs9fWv+7hlIz2scljSUZNyBOy9vM4kl3n+n7zwOJFCjwY2FX0y9x6i/pMM/7
cHnXaS5X9MWznrpQy8G3aPN0Aj5hgcm5HXLokJpS17jARm0XHHnoXtJRaqIt0ykDIX7+I6nvrIK6
2D10hBe1MG5URS0kThre4WqRTcbPs7vombqRWHwLi/Pwoq7CUZDsPpG9WIdNzieYXVfxoupTFoxg
BTdwpLTGpoJrBKKWfFcKjg69fEMyDc3Q9v0fyKcQQsD15W2Aa0NttIqhZpxJpaurp3WRLjhtjnkn
gGNQaF4IB7WNr3IADHoQknYqaCHz+jfkXsOm7H/73Jj73zmMWG3/w1R7EBDU9YHsOP/i+htXGkT0
u0+TqI9WkfJGGayGVyGvUYffm7Lf57+DDxnTht35Cw3iE2mKlH3u+ZLOS52kmo8rZ2JKuWyU10oD
B46EXp618m6WNhtUPZbgPaifDzvygZNWP7qHXqwTe9D8uHZG38zFDSWhn4/uDZW+G5jB83S1sbMr
6u2qxGcyVkDsjSRp5b1qUIqUWg03yyeJY0TSzMWcc2DPkQVCrtUK69r5Yy3sqG5hNxZAzFvOwDD1
ocBJp3izsWeuiL9P8NB19mONlm3dZS6q1iFltywL5Op979GT8sIRhoKI/CR5shzXKSUm/dkWS/7F
jrSK0Bvp3kWPjSgQJYrZSpojzvV7cp3B/jtM5a0Fm5apTAXSwIfP0Wlf/wdCWKoKXaoK40cVyrGy
9KRg7xb1C/cuPgUCMySZ++KP0eZ6cjNnsGhug/ohOsKgNtFL2N63Wl25ycXcz3gZG7ApOddH4v2D
znJfuymuxcEOTlIVFjfvbFTY9DGrKD8Ee33SRNjsti5C/kHYqWtZnVbA7NkoJsZudoNiy3yImuFa
ZziofV8QvD7SoC8IbQUS2LYdnfg0hbsGz/Mv96eTbUAO7Z59OQbDLcM76m9DcDpLxA4s46eaDi5l
PJ5LH1luMNsoxKfN13LNSdqp2miSMvi8D46hiOLyAzaHpM+rjcNy906pTc/C6nsXIsw8D4MRWGzJ
cnI5+DIcxLEbLaXiEjlvRYqlFT5EAKU69VAMGsKUMoyEwPjM9o9npSRKn3UljDLvU9V4htBLB4bC
DdriQiLYWdPYL4EJKIMlAnYgrsurjxcmCrOWL/s69VvfMmX+bynBHPVCCnJDjfzSeZTTzycAC9Xp
m7CoceIULf6wHZcCJRrB8wHqepgWdAy0KWCJdI/siS+DoRihgZKPw3+JehWFkOyc293Rvkyi4eR5
UxGaP10AJFXKbDZIv9KioUSiwe6MhUQxqouXX6f8ffs721rUYX/DdELHrao/cN/sxatNvatEj9eL
RkM/LlVYahhNoOLq77nIgFIajqnEo+y4yaJvcfv8d/IGHXzWqy7yLfEB+zY+guf0PpYJ/vMnUqg6
X/O42DDsPof5QarIfqI6+K25V9K67uZ5TfI6mxERihNemn2XnUKcGiM7P3vjxh5F5BOEmWF4sw8J
tPlvhbF36NQAPzRPU1vDPqDugKrkoupIJFfSxIrktBfW9r72Rfc68OkaEtqKnYASrlXQlm5Pj4gC
3jLoZJZfuJ+wDYmLc1h60LGhnON8sTis/3KK2dq/01jMVNgdnXY7YfidzuX5DIblogHkmlOOhUwC
USbtJUyPIRDwC5yv/6iVf0e0XI5I7aQk3RV4LHFZdav0VGx+ZRVHtGwSXlvCkcmig9UpNpLvKEHv
cwg1WZBjnyh2YDkhxrqN0S7Vcv5JhPLRnas+ICmxq4GvqoxHwE835mvw4hQYSbsJNki0tgX9t5S3
JoG1hq4QZTMwE/BA7Jg0drXH7UtGGsScVib/vSXAVuIRTQc5GLUOP44uA8YXzgfHhK+Uw6H8+U/n
KXsCzJkIGp7W7M6wyOBCHr866KN34Q71i+mUYBkTZqbao7OuA6go+yQw7JOBVCkOlN/u0UB2ZVM3
PSF4+qYvd+zElIuJ1UYWUwSbWkJPkD1pWQIS5nLFENYZbb+xHITMSfA//1ZQQnDodFQ72wgQTyrJ
pXptsI2mGA0JxrDVyAKdRD+7SYq/9mUpornfcpbT2MKwV6HC/y3XP77SJcG7Tum0LUkzm0ym44hg
9op5tEPNgiYuAGPvqoFVYDA+WZVicDRpHlb1bZJ9rRwoLFXdv3HX2Vvbx/iCKQyBjfv7hNwVKnea
60pMdIZkS4BdyT4W+pWuebasEsjUCgpwoOj9ticIV4r6tj+iZbxGZ/Ft7iXCQrE5GLcRyer9wfQv
i9DxYh48L5j11dmDywBBTd6a+xMPRTY6ReQod1mK7eFa+wcbV5QzS5f9u0UDOBnBmKuD2b76Fmns
agJ9L98yp98/eViNUqvT+BZ2kMjcW8FrgwjBvQ4iZCpw8W1/zFKdqzCkKNpnCOmIf0j+4OlP12ky
E+ePlqsjqmnY0N2OfzAADS1hIFW2HvrHfaoSB6/gFHCFKF3cJS4sQxDgv2denMss3BHrRMSilR+w
pDrniucqypsrdiNRzXz26xvD6qxKbZIG3zUmXNa1rBZZ1cCjq+t31ElM5RhWACGwoid2lPnfWOAK
n3tNLhTGzsvg5chaeX55QVjv19TgU4ieU2OEKaITd9Ghkeu6fZ+kAl75CAuHEnmIZ8vvz6lpFS2D
kDf8JPM5IABxYe4+gphp7d3I2SXAntLcBvPA0M30kDQkieujis25OowbM67ThRzH81vV1PeCdA0P
fu9+J6iP+lH8yWZCUKGcpG956TT5VcTSbVwqrNjsj4suIuo9A6tfD00ty9X6Y6HsolNtAHlx5ym/
jvxDO2MNg6wpsiAV2MfHZ4aiJou/MXoAdI/R8BusrHP82rwMJwLxxdKEmMMirNh404kC6k+QAju7
j7DTPwccDwCbcp7Ibrvfqf3DFxJbdAOSDYIiCi9D07ktwU4/4Thruv0bdIyzGIeAhKASJO0cyJ/M
EBKccD9Kx0CXJZCD0pRxYqLA5OFm1OOJK1oVSfRPMjYXYW2JmPc4inlEG5PWHuCLphegxSYGgYs2
v0RXRVHVww2nmdsjy+R0UvemelULiRJoL12etbzgm6wVV69t5Ox61jh95At9WESE0QzrR3HbSpxf
w9hkLgp3BsJvsWq/uv+oBVwMb2PYoX9o6Sk2s8e5Q+KVRQ08hk6W4v6YS8baLYrYyuzzUuqwljnk
OICxMPfVe38Kzhk4c4DM3T+KIOGjPwSm4PLQe4Tfe5Yoe5Cr+PlEeYUv8df6BERLXJ5J0N3eudJU
DHJHLREljpTun60bwPLVGWmGSXvKdNTLQ1a9faTGwTSaETUZ1khslsJjzTGcVqyzJL7aAeYZG96p
iX/HDixXRLGe2b5/daRw1dAvH39LuNe0qJuAj1NaXAIPeWa5qvxKykRePagQ6SEz9Vl2UDMvwzRF
Wpr+9N7UV1doGwnCi7BoVyexNNWcWyz+UnvcAdMoJF4dyV7w1T+j8mvNQ0FJc/gZHXcrN8kv2RoS
xwQd7x7BBiP51oNiUIn5hxNjSlHlCC+SPROzYSssCCIMsf4ZWUHUyudPuJrNbAeWm5or5c6rq0KZ
BVANlcvm0H/t204gbpOI/yjTtrVQSgC+h9R2JFsQ7sY76d0tJRVu3HC3b6rQ9RZVTRWEAqiYF3eW
Q64iLcdN2EBqffO8Ph8hybh9b1Ne5qiKZus8A4XcwEfMZpq+BrR9B7IfKoY/ymAcicvi5/JysVZc
4ux2cjQWaBEDhsjceR6Uut/3JLg7Z+JH1af+0Qe36FcUJ1Dp9DVUH0Hu+/2yXGqDAEBoIQyRCdsZ
zg4pwP53eAntPNMvWhPbkPl0KXshlHmSoTsOqRq85qGlIZRmETBKcfUXeMzEWbUG02ePF1HSWgDM
IZ0KX4aeODTMOEQUmKvmxigiAuoDXbcWjzAL2PX2FwKNUPmEEW+05/EeG8dftbBJ5V7wqfLe5G3B
MLlsFz2dwIyygZTU4s4zJzUKLiQlcazVOWKoWMOhrda3QfoXTZshGviwLRFn/PSC8V2ji/kc+AOc
VBz3bSLXl6a9iU1zARrE9PDbi9FUqyjmw6QWep4ilDuZQoSdmfxd3uXwtjJTT80JbWMqlj0o09ST
BCgaXHqQufvi89CNm3yEsdVhCvnofUyvHVPKdLrqdAuz/06/9mODWwTMb1fB1a6QMfJaYp+YJNvk
UJQ7KE0ZJ58vxTkA0gvgKkSYG6thIJkKOWjlWh7BfKNKDNnBSGk8Flg4IJ1xE3lVGRjDSdcC3hiJ
2riFa3errTOk3QmIh1V02KE0I+W30XwYK6VQM8cTZqTynFDSHFBBvBcjkXs5F3bDLp7kC8gkG0Sq
gZPCPoWNYmomQb15ydHpOWsrOh4skyTB0Q9y9NEotO2R2tJxczVjBqXBze9Vo2K0UKaWkFReA3lR
KEXNS42OWYqY8GhCV1YqgNHCIKRrZVfPEgZv6riu8HMIT4u1VIaZESbGPsWwS+lcnGtFvnXHjcut
fkBlEW8La1ZX8FoPnjOOhPt/7RGGZGI2/rFt7VXVKoOBY9nKPdl8JAyWgvCVzTlHbZCoBgO+QiGZ
GCJcx5MOo139bm9FjEfvkEgnzrDkiTKk7dTl3JRFVNG1u5w/Q2gIo9e0Mlo0Fc5ERyuBMmtVOch9
lSzHWbcav1jTwrNHJ3j5CSvZWE0or9KydkwwZ0rPyK8rjpr63USifvWfMiXdeu5Rpma8fdcrkl/7
T//Mm5JJCgFLk3yn5SbuVGrF0mGt9Juh0hROsbCuR6jMfW/94ZqHpd/9Vy8kohGGRfHpk8aEmfhW
qTnsTawdMr/xWNHtKTSRXnMLT+VI2v97j0saTwkotOHbCVTz/mTP12Q35earXViRuWc58QdfZSfh
QVXVSS8RLD6EB2WRfeEJ+WoNA9ZfRnU78fjXMPz0dB0glQ7S8vCBWQDD09nS7gtDMBXXl2+pwu3i
yCm54Nw/moXLujVYE1P1pf3IBCiVB8TqI2Tik0rKr26gORNvDOt3fa8LFJml/rbicrSZ1fX3I1nF
l6On1YxkvUDc5V3fu99o/zmPRyWQGhhrmYnBxG82E6QTz5YPRZizVxr7EWyNtF73V/REa6/AvL5l
S4vDWpRjsBCskuxzQy5PKGZxaoc1ghVPm+zvuuenX59qGceFhDdKE3ZfiIumOO/aI9V5hylSm9eR
AzFDSuxGG98/nowC/ZSFppahIfdUGYDHjyj8zdOi18zNvVOGumXxGQcWBHqT3xNU2oqVflNiCwBg
ys737XEJarHV7Y0q+JxuyVpwtBRMW+08oeDvyFZRDIC85RZYb8perU3z28rsn0lH0Budea1xCSeo
BoBPWtsWtLeYu6o7RO7D4Myq8qPgUGsPUh/S9aq2zEfm9AEkWQFQPuRsDYTb4Ps22zi6p9Pb1SsU
TE2VS1ukKsInrPEcUwWTohftzz58emZvcDwaQ/ED7rQbjrK1zOvkpIfPuoYpStcXJpc+Ew49qY03
Udsrmhj9/Ld6KFhtTPpQQ/+KlNUxKzR1fEH4qYk79RzQ/xk2By7BhvagcqiTgzAZSwQxIea7xVxX
6ElVrGS44u+iuIc9a13dzY1IHdezVJDtEUcWgX+rehJ+6eVmmEnKg2RQ2uq755Jpstr4NrJObmbA
do1eQDS29dHgURT5Y6Bkr8JTGLb6w4mhtp0z5FAybOALMK9Tqie2uogQ9ZF7ckc1AsZQqR8wGoA+
s8U0+s38r6j2QG4QbohqqTAEH9JwM40mlebkvXkAfbmPu6X0lq9yPfu20O4PF346G/ZcegiNDk+8
tTAKw8BmVCcqVc1NudgvPQhOIISf1j9nIdeBlPIL+7V25+dLJXu9Ch/dFC5DoSkiRHshbeS2YDZZ
PNohrgRlZ9wfDPYTYoIQ0ozTh7T5yfQAbUc02DdqGUU3TPjGCtcG8xkuuKH+8RnGix86V4+rQdox
QrurbvxE7axBIdAPnOUXgHiNeqaKGGjX36ujmb+yaD6R1LMYW73haawNCsvDBxY4pEW+V7dG4j8H
KKENuyxlI7/GaXy7x7XqtV0Wr7EVjT8ldFA/H0LI4btHHyWzRp2PfdKzkK9oSXuNh/UMjtZkZXrI
lsWirhafMklWWHPjL/157YZMGOoydiyVW302oGVoNaRHePxP8yqpB3Wl9y0HUWLpKLDXbwreJKDV
v+CZE6xoYkGJK8FQlXTPNTT3lTAQ/k7G5oWQNKIoC+BRN3j5p9M4BOD672HAjvSQBZRg2hf4umIX
FIEPKRXpiJ3DhLJERcz0ilLXHdPJcSdiMs+VV/1xmBB4dsC9PYoHcUEnUQOqmAzHgdg5CC2xsw/B
r62XOEcbr3EmFhcx3rXIBp3YSu9iP3jgVqRm80nZsPntuy6XNZGaHAKZqtnykijdmaTmHuMLFeUC
+eAICZFcIoWGOUHNHHAGKNbf2LQJfKwW1FCZlwlj2b51ov6FkH9qrMdgnUd7TJ1PMHj7n0qIsiFh
3DywfhKAx42Lkma8uMjiqFFYjRQxk6oTLqGEL73Q9dq9KQek91FwQVmIPbgsC9lmaxK40zAzypeb
M7JvY3Ps7wKpXw2V1kaDuB4VyrwcrMnJCt+fLCHqlgOfgod2IJozyVkExIHyigovPQGSTL5X6EHN
NcMxo71pRtHnEImGAdZQsDVdkvgfN/OlJ5MkePRv1GhhSAqTB9ZZZMw4fPxfmtphX+C7IYDAdyJw
hzEKpr9XZjHLBKQgbq1D443YiA8BEFfnGjyY+r/9CyuRbjNiw+ntMK0Go3r7mZN+NeKHE42xxqjU
3rPdJV0xowfrvvADH6ghLX2r/lx22c5AL2d/Jp5mcof7v0p1w+VIn9sOa0jwkB/AEz4m65r1xHRH
l19M0/LDCXgwk1UqZ1QYDVwFRv6Cw5CA68HVoOA2oj6FFuqXmrI/jlqHQFPp8wOV7+5xNf/HiOYW
E3jzhhM+xXGj0P5IS6z/1IvgpWnLkdBCX+u9P6WYk18kjwKxCECmP9aXAauBPha8ljRky1gcT8Em
M3AkhXJA/Y6uUB91DSxapUgibtN0ZL+ntpPAGjYKG8WIDO9PW/GUS27gjBWk3cpvauA0EQTbkU1n
dq6E0mrhE0ZY30mleaJgiWPzmA9g2lCyW42ptV4wytVEf8oEoedpRKAXmrdC3VJLgnPyqeJLWrhT
RUTa1RRrQo0D8Sy1fiSbbozT1tC8JLwzDczt7M24PnMNeZh8E14PndVOBXHt8hKkrmXE3ai2Hjua
90Ylc35Pu3f8SNMAVi2NBj50PBi0cjz8ZjlTLf4VyhqDChTYczRUJ4J9jBR4N/gfjNWnWnbQI9m7
uvsHvmtECT5Ky/O020tUiTWkzD3ZTTTnqZqbncJPyXxKv2kq15TMmjmXx8HPMWtwOx1vmqrf+Ah8
yNZAIrLnNyD5RPOsA2G7u9Pl+AJpIv7GneCssVJHUgj+oneVeWhLr+s1L7pp2RHEi3lVC51uBvzV
nZzJQzvTcgBJH8Hf7IeuFtF7pqwSq7r8qDzitJz8MLuXMYj/pXT7d9JTHIKniSzJooXyUDaRutm/
KCf4RRUrpOcW+cxMV5MPSjANNS/o8p2V/hoE0DGKQUY2fQz6f4mMpjjoDN5oleD2cOqacot7yA35
JuHIs3Y66M+Bb4sPKdXE7UhBhzMtA9U2Vc444y6CzzzFibehVMiNNxPYxkiHYbe0JrULWj22iztY
ituPml5jqZRUDdtZiIHQqJWxWaMbtekvcfA8a+c2kcfvDRIhmcJ/mvckWyMg8tFVsubd/k4YJCCv
5fXSM3ggp/TUwVga58pXe0dAinUXJ62wfWiiErz3fe1JyXaBSu96C9yF4U06v+tuMeA99Zd/2VkX
fUd2Ytk3zMZbQ9UQxS71O341jEih4LMtdYqhXf1xaOWSRYlSGOX8dA4fXAlhy/eTBizHCPc9SVg1
TLCkkQlEsc5n01EqGWxog6Qn/FcGg5u58uFxyG3pXTs++Q6BrTEnOereIy2kkNuwdzeFMNIDP2um
RuO0JxyPjeT35yjxseynpqyf48y+omp1PEG4UC9pLegzt1i4nQHcU4w1F9jpUtX+/+ls9+Y6Yf/+
cODtmSzquMIjROblp+KmBD05/5Qohpc6QHJDgfIwdjxs7O+GxJN47SmCTLWRe8RKNo7nbMy4NOAl
NIyzIqxmGSNIsjvKTAvkDPBx6QV2Jsalw4Y+ogY4R+YFegvkH1DZEc7/edDYb3VO9HYm8S746uvI
2WUXBlQhW5Ewmw3tHHBxTyIttF7fL2JUFSTpT4l5/9LrnhViSPMK7uSSzodg5LZ1w5SPMWgsNQDU
uAgvtmLAmLzi7X7W2vOHV69Ot7JG0TUPm6k5ALXcLCst+bmBZAHAbkzogg/P/TSdHJ5eSjBfL7yS
BDQmlwn9PkuX6jlNPSyORD18kkW/poZNB2yafppegZnUiCAc7Kp1pN2AFkh1axGwZnaNMLrBmyvm
ffBaTImePV5cuHF1Se4URFLbbXEUsM3woNMY2Ur8TALw/jH7xL+57OsV8yhZmqBJT/dHG239bbs5
YwpLrIENhC2SRTCdDXdFQq32eUFouzTCxU2fEWIggnW+VTF+gleic5I20Wx/t7+jB14I8ff8OGNv
1FUXOrmyXC7KRq12vY4UNS7roNmisiiEof0ZMKy+tEeiZexBhRSVG3291tKzkcPZ6xCzdSPAbkzP
KM1ipoUajfhz9A50OD2kxNrTTT+vHPOWqxC2O5njx/c6JPr+cD1DjWhuzYzW/20EU2NQNlqz4v80
hlHWEvc92IadcrSE4ao+DhyGkOW2njcHh5US6zl00WbzpHsdKPk/VDlB23mjoirnXAjvxyoihYgW
CNZ14vFyF7ThgfTKJYs4lj5Up0t5ZzHtjWp8hNG86ef/GOSKgcHXjMRpTj/ISLLAzQVcJwqKPNfD
XskRCvAXrD1xTIShla5VZbfQURrQH2YV3RdySciU+sSsqwaPVD49SkfNwmM7BwBmsKGqYXwvX+at
pktoOrVEUwztSwunD1zEIH4eAyIjVK5R/qrcXN+QiamtfgptE5OMY0NoHl9ejjDAKitIiCr2+TZt
Tqh5dO0GsnLOQj3QXJ+6dsg77mJakQNVsmXSpg66wYUCb0SQUy/+hj2vTb9dqPMy8+shkcrrb3as
9OXLuaAz92a3bYMqn/hrJIf0IZ4QevBfRhJCT8uCRuk6rMLkedhJ2HiWAzuhzkVwSJOPCChAGH+q
FVUaEmp2jKCgwVZ8Y1PVS4tAa48GfO/9cfki2Z8oBC4QKkDnmHm8PNewbIhWVCOwHBsdtm0E/94/
lLOmgrULADTIAQ88xZGiL6PVAyGUmhw5VYdYDbmUy8iRrHcuLjwxsxDkUogSMgAfIY4omupeHjjj
5QtM5ZvIyxFgZeGjFGjBnMeMlcIsELXPTSN/KDdeg4yRvAeirAsq4LSJN7UbLyOs60HxBzQyS+HU
xVajK9t//FPo86ivjE4XcP3eAb3BUviDpb3qobRC+MG2gTG3zEEyZlbGAdcCsfPaoBtk5zxvKxIT
DiWGDkuruoivf2JXtjXwQ90FIRpkPpkPDN52ok98A8m/aVNlttPPiNJpfKluCEjXVtBAgct+Enc2
vKHCo5Ctnta7WuKpx1+fNOQKHW88VcwRg4zdgQHe6UzG6MqJMFUFEqOBOBJoZe6Tet+LCptDUz4V
Mw1vcAuaEhQeKsin9gApD6Dky4VFRDnkRDaAqpRL9hWx4mvBPQJB1/hbgI5ZtmA7LkrTktHkU+Ps
1tc5L5ahgTPeAyw2bctTrnz4f9dB2YnFbQbZjtl4PYFjN2DDgILC/PAvaAJcvRsaFsMxdIPxuvCg
JndnSxKxjpDLiDGUz6AClEagSdCwc8nT0/DOO/8vHQ1BDo5qgKvRJaNV2BCtSNGU9YIuCe0aAJ2u
hUWNbB1vuZMIBs4bXIl/erDpIc8IUhhuv8uEveN3QX7RhzyTAJqkyBScb7Pc3kW4k3g6XnKNf0nk
zkFeL3tdnqBmRyMx37qtSEB2gFxJlHTlFXRh9XHLiP8Gj67OscGDajTXpcA9zeOs7835ypJU2BmV
/chUHouYW1saZOzJ/hvYGGPeY7Nh5BU4aPN0DRwALC9Eoyj5S5HkKIAnpFua+UuDOyX0YxOjzeWM
Y2UDekowj94p/RR/MOxHncCBib77vK5NOj3+uFS/p1mZAT/dD9uu5CFwe7q4HWhpJSS/Z+JUclly
g97aOGrEAXj/YV+4x2GIQ1nG7V4r7GIyXjTUzim51KMTAorOgfYnE4ZLZZw9E4oGVxyvYW4xrYDs
hBPWVwI4r4VnjA6fFmuZOK+4kWdPiFnxIEaHaU81g6HqnTYPN41f/bWz1+kwcnKhbLytJrwyvM+s
5UytCxW7Rwn8MCXZvoVV+0TS0o+pR7E2kAP5MEMigDfc2VW/hvV+Ynkci8NkqIgi+4rNKlajnDFK
+qkBaypm7LwvCysv5UBf18yBC0NEzDQ5twqVdW4gYfpELJGbAuyb4E1Pkgqykkn6ukjsawWyIC4h
ghbSpR1Cw3muq+Vrh7h+lcpBqZ0Ew/TAQJT+eq/+UqZQ260Q/+IuGnujO36488XM1q0bvqGj5Vps
77agN1Wix6hd9TnJNrNUzFebWaAdr7Op4X1BUVVOcwFZBOkdp+yk/OP8Fwg9G7rWOmv9vbbWMO2Y
hfMaJIBtOK9RskXfLNvQhs84InnfEL+/vkAu5iCC6YZ7JjgbzvLTg0yHlcREqexTmrjQJDv1Pj4X
RYDiItu1lstfPcMiN+6TJ+woyqm2i+HP0YJTRt8GU4y/kDjjNuJj50S+6XEf5TzLlDxXiM1Kyj0n
FZploxgSg0Ic/U9jNfyV7jS/8NBuqpEcAVfiirS6VKHiyeElr8fUdUHkhFG+cGxttUzRnOhoRGS2
Ae5WIk9gpTZnzM4oK37ywNmf++NXrvgeSJaxkvlLCMXprxiHTZr86As51O2yqxdOmCsuk9aMJ3Vn
Ovn/FtFh6Iajryf8ymO8KftpyGCuyuXjSYLd8lYwXKNXRn9ix+30hHHsd6p/OofMyb1bAQy8tpc2
a7FcqmaxKorYTori56R5ZC97exlW3LmfagXJ9BXFdG4L9lHyWlX50IFa4ADsSrTRCiq+rf81K6T/
2cSMoWl1lTSxDTbEKDpYw8+A8VE9Tq2ztCYH9Oxis6w0vfvCzQ7vgu8TyDhHEU1Ya8Y3dfAQDIXT
vkIzON+eSd960y9vmj8Pqemcj459l8A4+MDiMMYIzT+ehFstgH6GkWAGYwWtEIP5NZd7h4S40BQb
a/8D42LmaWh+3dHjZoW3inz3SR8LVqv72+apr88/BOPjW8y14k8a56yKAt7uGz6DsRRkwS3Viz7l
MvqYd4xvaNXBcSWlNNViYaFPi9UkwzuEX7RLvDM7b5CdTlh84z+4AWRxMR72mIXPFnN7zd1JLFXi
32bR95xZxc0qEBXdvWL6BxeIk7SOcLk6v7mTFrNoa+rlCVxY0tW7D03Nma+CPfMxhWmFQuKi/HbA
lbM0j9l8K/mPs3H+KCdAEj3e+cMTqE4a6jMaj0ie3UrxuWI2VljZeIBY0L38Q6WYa6nj0bbWV38F
K92KdWbhudRSdcyzSDRYy5LY8AtS51+i5lLyM5h9kgXPIFozjPXL2MLVzL5QjjI9wK29RsXIOiLi
Z3+SaEz8A93opAfFq04oC7ejHH9UmSXNezxOCfbqn3xXOSXotkHeuBTlGtnpLinqDIS+5Zr/kEa7
hP4enWhicrDXV6J0vVdyVQZdy1FgzCTidNXUS391Qy9coiPhnrls3ZYH151eIT7MeVQR5x+4gGhO
m9CDWQNFbg2LDJV4+VA7yVNtmAVCNCbsaGe393sHpet4TPF6SUa+EbWfDIBXg2yvBcKYdaSQoCP/
pWcNxL12q7X7lh+mnxXfVTn5IsCkwhhMs83aI//oN0FLyYKR28ult2G4SfKDyIuGoogHSbiGJXQV
ObvAbwo64Wv3ZMZViGGWfGqUvmlwx36Rf6OCNJD/5qUxaPs+JAD4/JM8krMtsUuoL5fWFEkm/6Ay
49Rmzbi6/cQH47sHTT3yk3D1lYwGBctabqYm2RqYRcNM2TYLWDDlDz5ff6DFaZGBPbvYWPB0F0kx
kCq8Y1Ensifj7UN3mRLpGlqANAefCYE1dEJJmBExSAoMdYK3FoIpqTTut8J2xAr5781P5Nvnb+dc
WbF9ge8P0R5PigT2erFPf0Pm3eyDe4hPHweBOYhQdSIsHrzrmJlOz0F504gm2XR4nThk7pmQFZvi
ZwbYfKZsOvovWW0ydlMdTk2XvIRiVw9pY7kJsKnaqBXoPe28vLicPMc+AJ3yTR/4w6HXvcpJH9RG
wi/LwVhzYTJaQBT2Eb3csfJhgKxQ3FHWaWFoa6TBbTsJ/cc8smCPh9YuJ1w93ZkfZ+PrIoKysw5e
cnp2ZupBgoJx2HYg2nhKBG46ydWdPoMEVOb+QJfMKiQQh6UqwOGcwfQIlCvonHKyYHAAOlkKkVr1
C4avFb3eFgMmhfO1feXTGy3H3/YV5A46K2LWcsiiqOUX3VY7F4z+ip9G5oM2CdUX2+DFC7p2IhBv
QxfrLR9qc2Odfde7igSGwvt5m088oh0aLELWNhAHe2XzSw10bXiD3i7ifAURUuPlfiIFStKSRcgp
pSum+JtX947VIIR4gwFFRAefpnjr6MA2ISoUy8n0mlYC3DiFpBIJrA9+Rq+yWfrTRQ1x9LuvnE8e
E8tyB681qjFdvboULQJFi4zDFuqUUtii4+psRCrovYV1pxs5vx6RWJyfX+AU7H93OX1RV/6mfk20
hHCicEN/2GcNdq1wJn4BRcphB68ed7EoFC9s0ezETvtQvDPoiBjLgo4O1uyqhMSM1l1gJUPKSxN+
miDOdkaGA5ejH9z+7NwkmwWEdj3OLIPBkJngshJXOYjORe1Nl0qf7Ej8hwYhO1krbg+46HrJ5j4U
GxDeMQ7BwJhjoPTtSUrWTJ1L6TI993ZiWeu4g2ldjzURCk1MRdZH6npKlmLxKYEJKmJw3bd6ugyM
7hskB1hIElDuKLrTjciyx0wLN/OrgKsrzF886/WBl4yzz1ERgdblZtIOVkWYZFHCWAzwpq73fHp9
w8FB7Rm4EVg1Lm0qhzYkXJYxE7RBtnu3Ufk0RX9Bh4SrjQD+ZHuyrrj4Q+XoaONe62SvsHav5eEd
06QhkjQqWYkcTNLPzf+ehE6trvZyp0R1UeNY5QY1Tr/Ex165GHUoxZ2D7Dt0xXBJ/Jd7ZUZ61s6m
xkUF0Bql9jQkLaAqpAR58NTBFpwwG6wkXUx7+f2lsiGmPDAx74XU26ZvhVZ6eKfP80XhWtSu1BTN
4777uusjLVylkUL0DaSG0NF8S/4JE8vzuClijy+WdEzSXVMPrf/C+Mdx1zH9eJWYsCLuJVSIThgb
aSlyXn2QX53GwFiaHl4cEO1PLS0E8IIRfaT7OY/rdXBrqZy7ssNfKf/y+PVeAkYt4RhLdroIdC9S
KoZVNcptBR6PmoAcdGt/YYGFO0m/WrQqVfN3HsvWACGXpwXGhJIPCQ/VyyyDp/OEktaGX+8+TcRn
k0BMA0m90X0Opn3XGLIdy4zZvCyT3ei2gVXK5VKu2/YweTy0+FLqu1yoxkePX077QR9G2vET8PUb
zdrWstc9/mbp5W1Tk5vvCQG7j6McbjRhRJzzhSpP8PNxEhcy4JejFugDWIFdLmJON+tw3Nmz9u6p
avmFxNy6VOd8ITXVfKoAywZDEzZKbj8B6ZJxfv5/POc7f9uTLRJNrE48mDsvxpkNYol9xcaPhD+o
A0KQUPJru9BxeOf+gzNCj6TenL9QOT5gfugdRqbnxL7RC0DdYIZyvMBroIM8MblVE6FGCB7qwKjZ
OKNQ9ujbu8OIXKdTw5og0OzCpcA6qDE2gMTfIrBd6nr5YetgND0+tWIHDt84IOmlMpolBPwE7325
ui8osrcJCqQ153ZZ50XKIjPBBKBAYg+rVsUkkLtuycIbusueeHijH1G6KXinGXo8zyR+LeH6BKyY
/Aq2Lap9UvYR5xlWcRfdkhPFxtM+IFI4pEYaVwfQRzvW33RX9FTem1MlY22FbfrqN9TIXOG0vBzm
264ZDQUNL0TRKVVKG58BOMmO4eT0OCLlbaN1SDIyRRau5UOvWx8iK94YqLNSgC9PMizmsOoHWQ5d
wGXXeTM7gNaZzX91opKHtW8kNYmmsXt3QYHmS16MpPIe1XseV6eOmKNJ7j5irx/3qGkblX0CjaW2
UNzBR70jU9YVtj0kUvl5yJTlWzJ6MdmZ1WeU2XHGg6ADzE3cA39KNsT18JrtN+3AGbe3SIfdq6v8
tizQidSAsRBpffthvmXAfbMSY5ozOqZ2pW65ECIpEzUC9S8dzAMfHZkSSfHn2c8hMJwLksUTxy5D
L4fM5q+MJp5R239BpCkvRl1FQR7y4yzWWpQ/sITrw2J+49x0He5dkSa/tXgb4yjmmn9tSPG3x0nP
+0zpMAe1t3d0QLL/BPfPkrIU+quBkGL2NzVAvRrwN1w9Y7eDt1lUxONDlUEGaWS2eN8nPh35v5oP
j7Epe0/pzEyl7AQirlXldxhOak9GW+9NbvxjkC0DAOenU7mNi4msKErDHnjlMVM1+Q3I32L/QBYp
fY6fxD8xyc4eJL4GByXOyM65euyRzJDZxXsc+k+wO9dWNKn5EqUvdrX/z06pthukas1TeevKpwxN
bevze5rfeWFFPh3ByMIs3hq8g+91oLtFDC22ObjIiSJVPrDwilp/qDduDs7X6SKwnIpEDvKNG/8y
pr2II4sZqLW5qi9sl1KD2P2p8dp8TpG0IRWgXggREkjclpDqfdTK65JFoFtLH8K+BXQfwp8x91KM
8ZnirdxXU+55mHKyhlThihhC4NhV1/yCze990cksKt3409n+WOvT2LDLVvGPTicWnfZxmGmUFaGb
9UiITde9Wzr1IfR3DszT6KfXI4O7BwyWKCdBaYfgl1TRpRjW3cHXWywGdiHTbi+iRqc/jP+fIydl
eTvFbodlfrRrFWD8M05YZfpm8Ej79N1kbPJdsxakemafxxuTKMrwNxjU1RhFQ65hcXzMZuQKXOmc
6ndJLdgh9TtJP4a4obRgU8bnqqkozbTpS5TRvOIq5amx7fbMfjH5LF19tZAnyjexjoG3/SpRCcGK
CpjqZxSV3ZFt3SVTYDqcRmIaia/LZC1eDnNN3Uxp2DWQBzIkB7+1IOYnDdjXvRn87jnNeFQLtboj
L82fY1wKcZDrxmnQdWxwAXkOjXC1dHFShEBrnsxiGWFHlgm5NcqKYKBhr6f7j9ZQ6gNvFcf0neJk
QAVd+bmv7aQDGhwYTbyjBeB3Jg7zYKcah4OR/pOhI98+ILcYIefXD3wYhUPtMTUHJnuQ7B2geFU1
ZgHTnBQGo3KZ5rO8SsNDfyrtCcepkZJQV8KT9crWdzoUTPUh4VISPsjCwLG+rixnXW6+5Se0T9F/
cS9wnX32GH3HtrvLEHd0c7IeWnvGR/camOwgMdvF8L+qtUzHKKr3ZflqdyfaG+ZzNtziirtdUv3D
Mh7uA+C5oR2stHSlyh8C1xWeNWF44dbtH+Kt5sysRcsHDdB+cKRLvkXw7LWSh3ppfyCctQY2Avr4
XIPNHURls2Gyijy4gQyaaPNa8Kqm5DDd4Zb6T9fRmFBTVUgXrmtDWbzL6LfvfWuYhrlixF4kIGag
z1m3AG55Q7ddoAy3ey299BEwS8aJDkASuOVdQvonOV/U+X9hDa2Hn6cyYNVv4OvkuC2F27l83xzU
JUrjAEjxjxYodIyeRGDWXnkVv3wnMaMqlY2nzK9eef7lKFjeWsFuDz3iEmLsmEdpOH7SGKINXsbW
OGRammpMgcib2Kq2A9bRooVDCPcdgg2ywmPn5Nld5IfD6FXptV5e8sKy0q8x1+aV0wnCibuneVhT
lZ3vaTCok/Y34Gi1stj0NgS09lPG9vp1cjKsNHmvIblP7pGVNrPBbte/N6tb7LjlWoT3pKeD5vdk
Egrp/iOFkETXksC70+aNFYNcGXxY3ILFc1C/I1OkYEWMfFkJQzyZUnBtf6qgLe5HnlpiQxh0DjYk
IXDF3Hg1IUHPCJfNfNqx75/7g5VJ3hZsag9WTXXM9rjvETU35TMI8Ndx5ZJferxwvu1t6W+sLzaj
To1JUysbSwsXQVgWih9sT+lZQ5ItRIFoi9PBWB7RhjUqv306ECUME2HLg0xOsUndwVNkJrsD1Ht5
/qe+dnrcHvTqbJBtOEpu2W2mrXlrIncvzjvr3eWHWDwZBeUP6VMJUeZInEQ+1ClCli4AoAQHH8mW
YwgnQIKp9f+hv2FKiIj0MXETl3RM+qFK8P0Dz0KFYv+GkU6mIn6pRVKVYHqhEP/eTH0502CFDaJu
a7R61jgN1lfWKL++NrQBaao2/QPkYSS5HNzHrsBz9+rdCbPPbF4HuVz0Zqw6ZkrTBCafbb8iVs5m
6dH5zEEI4aNz4uxBM5Zyb20zqXmLkwtcLVAT7+pOpwC9SIMyR+XW1cFHzPW9FvsosQ4Vrrj0u/pk
LfneQe3t/1VO27gnkURx123VK6Jk1dESfQmLZOM3e0r2XGDujXJTcyGRsxyfC/0yh+IMt7zH8s3e
aZ+eG47EjuIgBJXgmrkpa4ra+tzlPgBq4wCw05x/Da1RkcvfMPkwDq4wmIFPVNsJCKM9SpNDyE0x
nh5OPJ2elrkMzqYypKQq3mQrrmNrcIOw5dWGv/jN8ogwkUJuPokp9PPu5HObfI/6R7ipaAAykXuE
YoEV2BPKlV1DcHX6TmpnqSvsPUo/TfwMtI5W/7gkldcWu+uZIK78OEE85BNW0QxWScFV3T2Dlyz6
tBacLiYWuBLpOgL80kXEpaoM+O+zKOXjlHNo45coAhuT1PGpTrKnjiI0Po8XQFDeVNpG0KPrkK44
wHg+WL5d0KrkHqs6j3nXIvYaM/OKZRwFuqxmqhCIHUziI2l7SZujK+qoL2e22V4CeFkNPteo6tcr
aIf+6+05eMflGLhJp9Mxhxx2043oszjTnKP/XKuFtqjvn++Gbej9AdrtxAl+E6TRblz9URpg15a0
wfd5aoc2L7zvuvv3FsUJv2MnmMlKRYz0XCK8BHTPeMkPQF08+w2AKIgtbS28/4WBA7X4DIRrKGMv
uqv/oErGspHlL8oQoQgMsP9nzRcDr9AGQP5UYfaa0RWrCvVKZnUnyfGzzsW8gPU/s9cNS0IaCrfM
JcAPTMA4qpXmKJIansmxNLqxX4NNP4+kWXPLcytzcKPionfXe+wi3VhbBk+KJTPPZ6NDwACaDPMR
7NJ3a4anHP4+hi+eCckwkOUcHd/X2fOqu2svj0WZLMyTKLq8sUbp6xXlR2MlgY1HvTxoVBCDavJh
7MQvJCZCShX6nszDfx/+xsFa+I/gilt13HSYmCkXqFNYkdNp8uhHJ7GOtqGAPHbJJfptnx2vPEX0
jraZpMbib/gio6tSwtTOob/2GK1NXL3xmffRuS/ODaBgXwuhIlVUFkdhlSd1Jvqco+qc9H0jc3EL
Q4nFwWBlMJYb0gG/BX4W5rQyMXbOBkYJwjoW+CQE3561mzO+DjAEQIUeXQvZGwot8p+Bk7BTnicY
ug1HxP484XBkWMurLGBbgbn1/CE8dkNeM+VrTvxvTZAyFtLeM8C2WreZEKRGBt3gyAYm1SIChz29
w5AWtHmV5neSjTyJB2ctPDw1ttONPOCvJWGUnDq0mYXkJ7+AifMX7Sa3Bi6C2UtrSjo2nwd2qtFF
kUwGy8Wjuxf9T0l6F4413OoW27xQ9MsOT6NWuDbgRJbaYJSgcddr/jV3Gk92x1HER5zpxeWMtPs/
hVQ+Eqk4LDkc8O1ZFulorFsKWCJJMcSIJ0NndWTMLo+jsW5G0SBJGtrT+DZ8mpuUVJ1RF8KDuLir
H4tMdRwQ+sIVIQ8qzr8F+Dj1S/ZhMTCMGPAOFERgd5n2sS8TBTOvw9Gf3rxMm9he+B6gkfVkIFd8
5a7UeNDdW9vTRX6md38n0cjgxezexztYPKYxeeoEW0ZIp8+O5p51tTpWQVa7aG7DqkTEpb+tihn/
NkBVLjDLB64l6cEg9SJHeoAwHeNsBGA4zArOGsT6q/3wG//DFi9zGzWojPQDDvmUNCKfg4gNTCpZ
/SItDg9GkwUmBqaF84ViSjOulwtx7p3OHGxwxVqHN9DjCR0OinrlTFj3uKy7F9fQfKnWi3TXBulw
ybd7y1JMnuIHci/lKKzwQ2CBCIUyzx7XAvJ+HmwOAbFTAHK6XSppTixGY8AxEEgl+/i6mcSLN+/u
gdYz2TsPnqW2Xyoevqz7VXo435a83ISETwx95TzW4eEkvAsz6LJpngKdQAtItEae/0sc0Ar4RCWi
2F2CLXIGFs0Dlz638tMLYy37CllL99nAABOvyajw9jexniEcBOC4bkWwk3ZG+TyMrBiG5OoZuVQB
x6ve2lbEurtg8Mc5ehBlrLzx7rGrH7gndblb14Yih7D63+DrrOGghoJUqTVTodMFy8LezVI91ojG
gWaJ7oz97czyuO0izrObFst2l05ciWVle47XcmoMtxLkcDkGpGqIHEgCQTbtLTOPh2oEhOXgSp3F
7uKyIJMNTp5ZeLsInuzWvg4oI12I0zpUh7SPV3x4746bBqU4h6GCPz4f8PYk5U+ttuypeOtmqCLw
UzA72GjJLR9w+YMEtIhVdzAzh0dxqux9Lqx/wWk1+0UTtaY5UtGnSUO3Imdcj8YkyWWd+UfM4f/u
QQxuF4CheKflXA+Y4KnF4kUjC7D+OO23I9OscLzyqHU9JV9tXE5e9sF0asNg305tkJzlQzOioGZd
tf0JvN7QdVe9V/90ysv057D7uZLnJxaR6UIK0A/h1HiW3Fd5P8cMnNiOFDx2tZv7VmAiVCIcb4aL
YTJulCIk4ipaQay+rwLWLudO1sFkcf2hjxEn1pafLKh3dx5MyIbJ61PzczT8ADXqJpsAOzOX1QeX
xI5yB9RO/+uBBXTLgJTKNpquC7X9Odyo3nhsiLbw2256a+x8qbfNCRahZ9we3xbw4srTjAXDUDrr
CyX7mD301WLtud8eCzZpM45g5n88Z00+iQhWf07Ny1xZCjIyAnYI3v5Wofug7X8j57U2CM3KqDHq
tMLB67eqvVbKmAecORtse2WOIoDfifhhUvbTDFQVkNfO0qNRU/MeafNQgA1VrZK/dH0MKZbDgQJ7
tAwJqHu7/DkZ/cQvMTOoBw3FzpT6U9gdK5IugSJz7udnRnBZDbI5KKqTuHqliFThvZgBsevn2kzE
S9Yhj7jUvBBooX1BSOhgMrX7ihrHBCeeX46bZyc9Qzp4UcecPmp1tu3lpWnoLbmNZX5+PJ7bfBXe
GuPciczW0EFxKa+9+7HoqC2eryOsYZLIjY9n0EMt9eH35N1w3teT1476WGQBt8jJGoKct73skQky
Dt1tR6DpTRYPVLJTHvMvAnA+SA8BFGY8sca3rdL8eRp40Zabh8Q2f6LU/KYB2OOEz+dGROtuntqw
qq3IKLqwufCxE+GK5DNttgzAsKiaJ5+xXIvD06+YRjQ7+VoAT6qKO0SEdFIYsosNt4jC4jKJT/2J
5RZkCKtIu9iNL7+7Z+gDEyD2HZNYAjOEoLMZR8ox/d77xjfTlJvgwg5oPpYb3DwSm52qamIWuVS7
xnb+Ws/CluauLQw0eObAToV3yGdz00sD/trDkt4EFWuUk8fbLtJL4my1H1rtm3NlJkX0Am1A972q
vSSDS/T61idw5RVHoMo5I7CFVk2cD+WmpIf63S6MUQToYc+g/kDokE4R1onKJnMXP/ln8+oiaImA
01VJy0VVojzRgAPSMYt99iKzBx8oO6i7L2IpXB8sREbL7Ps6LKwUlCocqYq/QeV8+qjBic+pGmN4
FFsquYY3J0rsBo8cf7GtpxIiTM4htw7C25NlKlgYhW/iAuU1buTSa4sEHp9pBUsN0quhfJVvw2gA
VX6nb+9brmCaS3Rr/nXgCaDnTAh1ue/wXYbof+O80HS+4LVh6+VKhtof6QBTJBlrpBAxsEMY2kDW
9BT+QDIPvaZZnT8Z+ZmqsZf9EsH08YOTr+8e7J+5K3LV7LM9dPu4MzuU2off0eaQZ7u+2aQ8tZgG
uzj5A70cyM4YVUEJmun7vA3APvh5s9uwfcHKAJY1Lm6H6OpB0iiDnITvj5jWYozCbDHyPdVo3Udi
FwRRGQOUssS/2PSm1YAsuNpiJAF0j73hwZmfZ1WuWVb+bPyVJMRugmQKAN7e8CwUHlPgbIvo5+ye
yluRGiIQSIJd2840TXWUa4N05ZS31CeVc0RHlrATzG15+j0458qKjgJO58U+empwQOf+afXBvoCC
Pojmf+TTSdiG2WyWpxcnyVn1eJcz1oItE5QD9s01KiHI64Il94lbkJtjhAIHbkZ4yJ5T2r/GNVjF
WzGbRhlD4x5DnkifllzOkrCAmbd9apYrC0ZaQTKmrqFTJu8QVJ9jFkENQRqIChK+UKD3ZD46kNo5
6tKHILAm/jCymSF6xjelecrJNwfjdiHILY2A2ibOfe+8Xu5GGx5bFVNuhtPYMJiHdCXzI9govYU3
Ajg9gQcGupDzJkZknVeBoVM6FFopNcdB4KSQM0j+uZNArAsJglRDh0+jhiumiHM6pnzEkU+uYmMW
NV2AuXybH49Xr6S0Z353LrqpsMmi3OR5rFhCoHvfsOUMlyOiYjoRpcNnz3gzIcy0f7fWBg4XM4Yg
S+l7igwV1Pz6sRw9bKrC1lXGYgsFe5D0XIzZ6WzldctRhVVcotoxuvjPOvFM7+E/cDWPhtmHOO0w
PLmMcOZworakF1462j4ttxutys88H+ZEuRry9l/nj2obb416rn8PEN+zxZM3GskN7vG1o5o1/MLu
3GSAcug34f9DbZonPmdgaVOXvK8/xqiJ0XCWoeFmqEzlUWcSNgxVi+6HsdHWUrAmwbyqXAkuHxYq
KpW7ooCIFhEnAzsTLY/iwUlxvDR0ukSKQuVjgTyzTn7cSOHzTA+18oVqn0DRtKDISGupzS+mum9Y
KriBkAFDBSKGrkm5+YguMdBsWhoZ4J3Ecyke5xMhQh8SlWGISMlY2z0pa5rbA/bEBOpka3mVdRGG
Fz8mEcebUL+WxJyUK9IugKObCVGo6TUR1XIQCL5/kVds+QxUqw994vf3lGfsZq9hzl7nx0QzJbhp
p6+hPqzs4SBbCCvnjJHpI2XNIs8v8byNPEruVRI5bahdFYclL5ZuoSmY13kYz5IwPogPgRvVfU70
4bBRSKrblinq18TwikHTGHuWaK95TXcJhlqAc7PMcrB/lutnnZewHFQ2cLk/nLVcUzWq2e302ePr
Qer/flFLKaZCvZKB+GCPCJ0dRrpwwyWr9/HFBgJHWJWWO810S9kdVOYbLOax8I/UKf9D7oIr9UBP
6p0k4XUTW7bn8pVksFH/Rw2401k/n2p/WnptQPb+84wvo29wGA1ZPUbkdeo5GP/k0WKbdsPuHDth
o/fBAGJS97Zx1K6z7wo86FCXCESjSWPw0tHUNjbMVURHlpWSNYb+G+PE7+KQVok2pQpDiAEjJi5c
N6F5h8MtQPcr43AY+TrT6UWY60364gSUwSolPcs/FC0DpaDlLwtKthzg4MZpLWgC8Fm/zo0a1YPG
tkkz4/QE+MtqLP0oTCHNXvGBpZcalAQKhhPd8wu29BW157iJqekgAcpIx/64Ec0MKRFibRuR8c6f
60FpFlsXgI5O3LQwKJ7bA5oXxk5A6ISd2cuUMT86G5zW7F92zwvC3ZK1aqFrneGQcC2jvXsEHM38
Emi/MsZhOOdxTnVfRqjGoXPNRiJ19selqEBdDQKLVeIKcT7r7jmwufycB1r5aOiVw0mC01Zit2Cz
e2Qr/0t8iC+yOmeUqP8bjaGpGgBg55Qt9M6ve9Uo2ZwhzhhIujC7j1nBer2e2y0rkKz85SHINKud
6KPyp9c99CwnI0SicsbhXyZRyxeg6pk0DkRZmPiwVS60g4OuF5H2r9bUlTdgCSgIoOZRbZq91o1M
i/mIAbT3zVqCgECcMy8CCQaF/OubVxDpLcE7wVF8c5eWkujogFsiKtZP2AiT0+AbVc6tpZxrcEhu
qJIe5Ju2GojHlFUrqs6RsO+4rNvs72FK0GSSIxCc6zQJ5J7T+EIugzsR4q4yZ3DcVhSHgd+U0dIH
QVY5LTfxBhoVv2HjvrWZQtr/iyuJmZ8EbBZykER4GE2NfaW37kisPWdqp6Z2LPruZ2FcHJehF2Ml
Rb6ymIEtKrqtfxfXZwRFtGaCBJqzkkwQgyhXRDou+ExwVAKFVQ+SoltKk3lgpw5U3CyKZhvUkKiT
YCrtrZKho5d3BBobnbGsctnitKmfRGit0XqKHfPQLxtSSLdKIt/sanQyvO8gKIyMItn+qQva4tJJ
6Pbm+iN6w950irHD55er+x25/5iPeh2x0lRL5hOylHVoToyYCxiP27mis0PO9lD0Szj+ZTYK2GcO
9v68DNiHi8m+vg8iKgcjcCffCvKSdzCVSjn5qtg1XWwXiVRut4oLkSlBtLnRnspjB8XI3KAu2s+/
PtQHfLyzoq0pWSrQByOz9+jV4zOFlEXGjpj+xjPoV+fQNlsdE6jLkICbPCdN+fl8PUVEdq8/7D8J
gdM22bJS1M92bnIn50cQHTdfZ/PkePf76woDdXnMC1RpUhVfdMON0w9Af73vRqSlD/Un6g8XYztJ
IB0g14bLsWp2zcZ50SX3hmiEOyAJ8ZEJZetvUAk9o9c0ylKlpmVKkHmL43bsRm2n1mMiw8ZCzDIR
93J840nd4b2cTSQc9rh1rAiiN3HhvVDPo71qAbV9bp0AP7bK0DNu0itD3oOSO+zCQTeqgQehRBHm
rvjuiyF7zMVd59JC3D3S8TVILAoxags1ax6LlrtQeTg2GVzfdzuHyguWrd80d/hIpmaF92wb6ZCj
WYFNGBBuTtIrfTWS0A34vsggTCKOrW7ec4DhorO4Y/2AiKGsTXU7JO6YyjBH1R4vcr6ZdUvB3cJz
+vJz5QxJAwwkD5kTRTLSW6VWHeE7HglMtbq2BMVjrKKzgHYfTvk9jBqfe8hYHqX6M78PlnMq+rpI
jjZg/q+xZEHneHHrECWsvKHW/j6ABvxlB1GXv8fGVzFV2q/tOeRMJJHzuvL0WyMyLbQTz55t7HRl
M9DKpY+6vz0KPNBmvDomKfueNHcLJVhSeQjI/iv6vVkGx3pvJCLxHkwD4jJ6xeYfOGhiwWnYRaRP
RSV6Ktj41Nag1BTD8d0msJaKObnrusYxXFfQuqqyBKBN6v6M1UlM67zcpafe5EMyuEfoSjIiynDL
QETkX6pLvwGKld+26dGoRYZUyQDuc77ZRYaKINRKbNK7kKFLdrmlgIRUFCmK+eKJyulHJ8XzY1Fm
04sq+7PcFaxrF4nZlz6sC/0tKpeBCESRZX8R40R2KPZb59hWOG9zus29l5n8pBtIomgioYDt98pn
9t11+8HfW0+v/ajBt/p4zJewkeEV7PR1HuaA0tZDo+yisQ0WVwmHlGRzeieBA674rFnJM18LbxvZ
mcJB+wDkpxT6xq973Rucg914+Pa/BJTGflDFThxyCG9m2pHVjYJjJ/J2sQTN8Y4SwYpnrf/LOaWG
TKdJm3AcURS6Z1M9g5x4l61IMongsix0Y2EMs8IMKU2gCPhNx8tT1kcW4oislSasz9+VtmAZXJoh
8M2jd4G/7PO3zXa0zB5VUtUiDeH3q1Th1QLxLctEOgzdoTQGg6876rBRBZsTpH3/OXMbFRhdgeoM
J2R7r6PM5ZC6PFY7mDTGeGGRXA43prGJJEtgzdtKstTtAtV6+FY2c0VA6/bbiVu9CrPv0mWG1kGj
bA9xkC5Bzd4u8I0wjUYHFHQbR4Wstkws8j0IMBan/wHfIVtMHbiYtsyS+YTZKdKb35LpKwP6jZLO
Ya97L/BsQ+Iu0YCpYf4N4OFhQ08Ac248486CKbBVRLWzr1RMGlWzGKloCOlcnFavYPvumkC4ujG6
T0MO1TC4O7/BZrLwik37AHpkZwBuxsG96PQiR8h44hwW8JC8f7YxDI/eaWSMktxjNbgu/lReuaPd
M3wn11q/XZr+AXGhN7eGsgEMHGRoYUj9LZmnIycgVvfY2AANg9235/rkX/Hglmbp4QWIlbZMzKzI
JWfyhm3c7RW/WCzms/27K4rH7lfT+96qzZAc65rk1CS9wqvXrz37LgFrp1EQLIaRWcQhx3pC+AYs
z05XB9XsP5hg46+tUgrRZMAe7dg1E901C/4qjfAh7oGFi754jh0lB6r/pnv0gM++vxs6vRqEn6Sc
dGhbr5CwCRjp3Y1E/BSodib6sG1BjxY+wRYgqGmZSwt5EZch5ZzCfToUQk+l9gXsWiSYtY0yPNXf
PxhE1DkbHCqU7s/bD78SDgi4lI+bEUQmJTX+SF3wJhc7cmWkoFH1fJGrOffMoB2wilVT6Z1C2+Xn
69WEyrFaD2gDNTtS+xyUlXp08RmPEDpwOXDCpGkGTBr0N+tii+aLSTkJAfwifC4IOogaY3OZKQcF
y/qtGlNnjIbpE7zob9QLQHNK3mtMyjPxiG0LO+ElYxa7JFu75TYzJuBF6A/OILIyJ8PcMhxf45tr
QcAZ8txZ4IfHjYxaDAIGuEAelSDnqc2WNMVUhFtt7IHVu441mWP+Khp3QoOjKJ4hQp4LGry2sE1I
ZBKMVovarM13Y8d0/eWIj5q+PjOTZv3AI4Rhvru8tt8mlh3EItQ2KpIsVPMkhOq8Krbb749tW5t6
fzF5P4FoHnOH/p1IOMgWya2Pfjzd93NcClmUcRcvOWLjhdvbaiMxvj6D5jue9jVRIJeZjFobPsB7
/UWIHRBPQhIIunMzpuN2huZ3Bdd6Fl1/kIwnXLOuQhxJCbGNj4eAxPk1/3JMfyjDwTBctPyaEsFI
kjisrfUqrJKrHYbA21g5J2vNqkT+/N8OKRZk/CzSWRn/SPxJAr9cS82Ov224YhPwAOvNEMbVw3Pl
CmuI612Uue/PqV0+Y5w/7zv7zu1mCJ2itpbYJtvX0rRTpK8PdFUtG2CPWzC1RbBWMXvYazXw9I7h
27vuUfZ7M4BmvcfAz7YiGdf1eJK8ExgtByMJsizWHm6nU3rMKNaNw1QqPcofWoJb+vwLeXXeVTcr
yasqGViegeygBb8BoJyBykecnCyGiAcHCrWJvdELXDcDZc0x1O2Ls2u9sfFjM6FVNgmrq/3W0Lg1
qpf8juQmD28sxhGwkd20ykKVnlEsNGzAYORT6FkA39i7sKN8MAKmGD5dcrytHD9p8Hi9Wj94XJ+X
qO7QTpLbT1fI9DFI+AS2W63JqMHLRIZOUw6QfM9B6w6WCdYczzr/vw/pIu64v60IX6bfaecOAdL2
Rq/1lokfZRzqWUuxxj9jpHE72K2z7joUE0ZFsRQW0lX0tZNhsCG8b/sDRCf8b7LXtrzm0GwyMucF
xBvvlCp7rVowioolRx6k3F2IigNfzqh7HC2bQDUWOpzUZgSg7szVgC9j4Ym5qgB7AfpJTsKGMPJ+
axdUp5lgSseHXK9ucrwwmPHWPSUr4yN4syaqGEy9YV+g3DBGYTL2vr6HY7nBgg4EhyQnL0TlTFh5
0EmUl4ZyYoTEQGxx3E+J9aGUyDmwl36gx2EgY7nPK1cH9Pu85MufqOq2mPfJ3zKcnCVsCC0NQADE
nFBO/JZ+dD/U5WBChmn5oE6a3ijwK4szurZoY8wlhKTMPniTP22TN+EWRmJ+Ir+2gTW+mGiShj+y
cfFfg2SccHrLINpKaxuvmNTyr3ZrMejkB9CcfDHgYzoWDUfqbZEHThoCgvLZtDnOdUzDkOu3CrlV
qFM0GK8OSCKBEcrH6Yikqr9SmvqR0QR3xbkGx1TAnvXsgx5eFId8pY1KP7pe7iNvTmPLy6hikEfy
JnmJsnS+TXS9RIY5CZtFwPxL9TQIf8VRxLly4tG+KdQfwNqr/PBJqFr4cGauKmbcHnFkl1Fm778h
oKeCAVXIg5rhBez71YewbmSlDjzwy2mxjYCIQKsBduohxxeczXxvDsTtLiGHgxrKxrBNrfQSg+E8
HjmBsETG/aPdI+t4pktRS65KSdGKq5zJ7GwqukqZu3/jJ5c4H1ku3nbt4n2uvkN6b8mCUiPM+hfN
DW9PYEqGHP7Fgz6k6UBP3DkCy3O+odaWQXu9hizsen7HoIYCLppp15ltZBNfXSFA27R/vg2dyIpc
pub55XGKVpy3XN27CAm2iowcpIOOH1yGl/2BfRGtoHrtoExef1SluLEsrGvteYxZpbumz50GYJ96
8ERX1KgOaMlcsW1x1YPaP7K1jgHb+Vvgc0nqIfuJ7NA88VV4QQF8xd3eLIhb3uPa6g7vF27QFkHh
Qo2FHMAieFD7jfsxdqpKPg4m9rl4D+CAGfBYdEkFQiIscZ9XIGTk9Ivu+xhTRipvd+yQKncKog0S
t3AFRsmCMAPpuevBngyXelDB9Hi/qOylDr4Dooy+X5+StK8VqhzMKsJzj2CuSOxV3WOLKP0TEGt2
RKlFXKYSDIgfQj9rMWBFql3dwbErRVZ1f4FenYiVIodXBfM/pWK18kMCQe5YtSPYAqOiE6/2hGnm
pHe/d54X/WXPgj0XxYewyFE4pw/5iK47bSRuei33wV22O5KZfs1j1hathLaduvr0HEbitinbwhBw
FfBdyW7GB6XcGRizVV9UKRzF123Wdi8qrdrEXyg6WKDdmHctxLV4yj2eoDtjZj+JjkeTcjFp6KVe
UiOxJqhbJiYMsuWiNqHkyBDS+XGfT1PzlnJJDycNxCGk6VD2D7E3e76pTk2lreuCPGlez1kklS8a
GwFFsj7htW3r0QWOYGAUJ96M4WKf1C6ehYFfSPoNSC+yfRRsO0b0Ur+EEWTOiobG2ejgtL6qk2T+
zWydujq2b3Chogu0CjHGMeWVV+x3pxtPkc6as1TwRkYaa49ajfmnV9eXhWSFQ2SNSAQrJ77uyA/l
SMdlqrJYTHUuZA6ve4TFmDd3e9fIz4Te1Xig/jFOODAqI3+M3cPgiG/gbRGRda+/mxmZ2r6T7LSt
ViFRvspEgbnXcWOtAX2EZvUtQfoi6D+9WTICTt54oiXJ8yxZpx7qWFXV8oJjE9zk45Din0huxRC/
c40wt8CMSouvAVW+S1pRVt32FwXIbiMwnNWjLWDwJJ/UPQJblI76WkOe5Pydf7VVhg6KsOoClcoS
7xY/jWKhI7cQFgZvCHJKX19kCnkdReZQma3jXitqXwXKEQNAovPdbpZXJqprJZkByd7Vmc6M3mVA
mL+2m1is7gdPvcqST0DHquvH0l7i5tY2BOaJx8ff8KitXadQnZMBqTGaqlA4xGiJMZPaDPvJ1GMe
vTmnMdOuykTg4Yaf9nNkVzZz16Q1baaOTn/xHTVpmtyCVRHJkKrcpUibWeyEtnj54+3l8xxevTu3
TExgi93ctracrHyCtOKpQpTYGCSCvS456YeTlbxeX04sqEczjso7hSwzIRLhWRLQPdvWic231Rwf
OvuwuJ+70XMz/g1TBp5CJ6C5rLguNVTrwN/PyioWo2/G0U3/oQ+ZHe8DjZSj8WUcK0wrKrq0fcPc
Dru7SBJmWQ+tmqmH5SD5YRs6FkwGe4Ccp7SvVA0xkJbavHXL3WN22PSgrFgLrc84SLdfe+lzZLQK
zqGqKfWWw3ZjdRjoJVL2r8HfnTENlJVzJoes5uNnGNuJAWz7tl7OYlWDR63UjpOB29SpRbIVvHWC
qEfWeApO5qmSGTt2Gez83XV13sdT0D3FV6y+7OKZMlaq7r+1No7V/HiChpvQpfp7eVkp3jMRyMuB
OO4BkOthYn7w8EqVdVdW+WTNrS/6BWAHAlD54aOxqvEiWFkm2aQKFh44heWDiV/yTW3m5Sfncy1q
YcMwr1Jr6dsn0VrTr720eRGRVYCb50Apfm4oEdjyaRGw6tn3pkQ1oua0PZSsjBco7p0XzCT6czFL
ptg0SaviDXAG3fpALin+bQNGXYDigZwEL38/vUmXAwDRfxnrZtmrcLBeYFef4vKkqkH3XQI0O0Ez
RvdZuDs+9ZEKN232dIiFtCynoAer/1i4lZfvpsGBHbLyP+4v5W1HXW4YXY3tzmRTdbafn2sOWGKr
Dj+YmUdjUWHwdGEX7yEy9xp6aWY3TnsaHlGVEdgsSWrTZBijRubizSjHMHsXTWyzT/QlClsdyRay
k/wuWMMDCv2EG5oVTnhh8b4PKAaOboGLxilSCY/tDsfubrv0dy7QHCJu0FEv5XaASSpURHHeH7or
JIASv4bnyoIVMmB4PupOBctBK+cFUjXUvSOBwBHyv3RR2icp20VM8Vk263sPU3cLatG+rQPv3lGK
6lGS9FKYbjZV2hI1zVqUvocj6u6w5DY0NeytSa+a5NchQetAxGgcHA90n8SdCqzr8aFP4ZDzJBxs
QSvBTgVUMjx8dP4l7QeDKpv81qHdtbTxFAUuBmwlTei5Ftd2axUfjgs3wu/bC6IhvUT2sY5ok5X5
y6iaouiOxN0OtWze+xWAhgyo9cVPvKX3VuWGfmN1aNRnH07SaOUuRRxCSV/nm6qJ53dGmnHDUEvm
ipj9KUxEpzI36beloASP+QCQmApL9u2cf3p1DFBM+kR9GTeDLabwYYlrVbLORNzd3p8Vc1QkEiyS
xcldAKNv6aGA85aPglibCERpRq7qo5WV4rFEkdrFg+S+jyGY6Gby2XfCx5Pe2VzAb5auKatup1xM
lg52qUTsbJRaYjELyUfpKBEZgB3aXxYgyRZtdm6PcW2puCrnPLvXHthsM5UZ3N0zTw2uC6/UOkA5
AhjuGbQu/rtdq3yQuhblis8ZJ3a8KSyqP37yPgOpRGQKYd6vz5GrD5cdyQIUc/nAD95AyMHComOj
sxV+guz6jsv0WQrfqlNA6UgGVYEj0wtoi677ylQi7eyQ5Z+PnW1l5/++J447tp17Ju5nJFsl189U
jlasL2i8h/mScJoi7UwSinK0nVlaUiCPqFist5FFotd96pUuqLwHVv04lMeArWLni+aW9MZsCf1Y
RFClrO1ul0+s+ArM2sIdTythj3oLmZJADY2OzqZUXMt+U5WwcK4mmiR7yBwzqoh/pCLISkT0IPZE
zxGawZgOY8MTDDEOrfMN1YLoDo7N02ddH55Mcrh2YAg1IwLj/BAmeEbF+FZPG26q4hUiCCAE5znF
1qFnUDHAtLGNLqkUHIi/sJP+ynNePbX9WDGxTJB9wiBAW/O4OEc+YjMCPnHylyADI3k9fKVmTJGx
YNtZyxKacomleL7MqcTQ0yKVFh7kDSpBRjAXZi8BIRdhUzjAqf0brxRZDjkgxcDhqNnQJcHY7DO+
7xRjHbNhTxo5I0VEEzJL7/acPbJu4n4HUiDP+Lcjl9I1Q6vquw4mfiKxXwWWJ7PhYcs9pKbo3J7/
UcORazbjsdGD+c85Yd0tobD4SYDKzQcW3hK6DJNXo0+uEjIMfSX6ebIidvNsE/pt2n6kOLILw6vi
7RFsD/a+S+1+C1nYhIplNiCNKs2u37Gd8+/Ekc1VnwuS+jWj1IElHwn4obuM7IugE0TBAJ0PuFLz
bz522mC0LsoMMZFRqwvDAQ1CIQeBk9v4xXhNXN3RryuO6MhEijD6CnG3+WOAt4KKh7yc+miXuska
AffBZ6Tb6zJBd8ngM3fB9akt2AbxcBVnMEPNGnsUrlXuDj2AhA8sgerApy8O9NjYAKkT8uYI8IgS
OMuv3YhY0+7Bl+xcBNAMU7hjEztY74fNyLY9VYWddqsagU4wemg6z9n/vcCXq9LhWwCIS6E3Fq19
r2nRntoi+d0P2KaiI8ZGnSMiYmv5fYaSJ5eHSYyEe5tgKHksE1KH+zM2M2yeRwNQPiYulccE3m+Z
xeu/j44133MNpRY4RGM37sIlPl0rSvGRDG0s7nNOQhY3Uq3TwKqX2B7OoySSlhHUktCppjGmcyoe
a6tXgzFjoUnBGJyUh60kjsJd1uln901aqo83ypAoLqCmUQsfKErVXsx+XaFU7vxXIVXFmJ0k5yiC
UmqT0ewx1OBmpyTDGxcWrDuTpQjwbZ3gFt4MXZBm7i/xj7RVF52Ab51qlUG6i2q65YuJTLg7A77c
wJwRCKroiB+wPKZVTHI0dgrvD6sX8gDvQN7sjU1W5nt84c/nTXS81+ZZMIKLGPzZtWjUD264qeJ6
ln12VgA46kNHTh8kz2gFiqZTVFHFBjUuQtqLUOGkFS4yN2LCKHMolUeko2VFVzH/lIQXTXCzB7N4
+KJ9EFnO/6Ut4S7pYmPLZHkb1J4SpijcFKy5060soY1+ozNA5oqXHVNnE2Wlrr8ea494yuDQuvra
MFdQ86OFe0ykYM4XNFii+4WlMUq5Y0mZZlvtw2s6OhS9Tq9RIReiy/6LzugKqVm4jdxbOOMnSgeT
TkNYNhbO+2I5sGQOzQTODm4Oyz72TonaQbaJUJhEfLbr//086rfoBkR/1NO7r2184mwcmv9oH02S
j+fnZq31N+3vuxAhNujDI9Td9HEEUerKMbDmHYMd/SwZ1AlvsUzFoD4aYChPd3kvV7T69Y6BVrNE
6gIpe86v02R9JbrbzFMMFpglzHORwGf3hrACwaNU3MrWd23hCyT8cXX4z/MLuupl1ZK3CQLbGxNJ
uC317ShP/jbDOie1cOgNVjTsDIVY5l1vZYI+SSnY5B8V2pTuldp5PDiMoa/ylg8+EXKlhkMY8OV+
bWV+PeKaYjjBSnjE/xNejMZDtcxlw+TD0ezM3z539I6mCMSOY+JE2gaoWFQeZhLAj7i9g/APZhSi
5qhTnKnkfMyfp+eqs9XZ9jU6svxcBBpjuhPVpz1HgKUdc9tIh27w7ttYBMtgdGKuutfhHJfWN+RM
njnndH2/n7ehIr6h6W4tUL90TBnyDBvKyETHez3AwjJJQTxRk7wo7iwi9q7LkYSD81S879iU3ZJJ
yetx2CQdyUJD9cp9+kpT0MndyfgzxeRZQSEY5CEgJYYjmZ7xWsgd1Pu/Of3AUCdKwna9I0Z5Q7x6
1/nUrBwk5CCDwIJXQG73OA45rUb/JpK/Ll/NNPN8ZjHhQiE8HZ5NwCdhRmSPSp7aAO4yGJbJAyBF
oLa4OZP96IRl5jBEj5Lgw/4XFh2M/QdkyEvq16UOUMj4V9RWoQY6twFsq+GmbmKJUcGm4EfG69zY
NarGcPzmUnNohQ7sp8lzn8RnciEyvdShVOxpGiVCpgkUdcGeaD01MQZFqliobID/bi8NrrIsvT9v
JZB4+4C9dhs4m6mMCJGaag+RGZFAt1A5LmCqY7r5Z3x6Muz+uD/+cXTU54k6Hs7CDS3qJ15vjuZ0
3IjmG1Uy+lr7fy8LsTWu+6CpISwiJcCirk6LiRdz1rrJ+XBV6TeJ+hEHGC60MW6Qo1a7xOAIjN5t
td5/yMlpweirtar62TV7NvWXCbXull1K0aA+N1j6MCZqtW1dufAJVR+dCCs/1gy7mdRzkbTZdRQT
AGgR1wcW1xyiDdnSl7acstp6vX/EJVN5kSNlsMqcfOteXw6MGksTfMibPJ8NfGoKDvN13UIcRpL9
ob9NLLRjeSMcunRxdDC8cm8ul1gO6BTJxPfGFk/i3n38aiayivZaLomcvfg4uRIX5YeWqhAX8mb6
VHqyZ9ka4L4YhuIXmvYUP2uH1s/5OfLRMTqmHe5WlDaWgWK4RRqM9iL4CesMXxHsUp1DK9XAZv2R
+BsLDff4aGDdruTivDfJtQwZR/UsZTqByV1MWOTa2dVgDiJd56RCHUavgmwN1N/5UVGFVDnVCIqR
8H2scrSHUUuBjP6fOO0zyk51MJ7QN1KE0YZv1SzerpcHKIZS9cU+cDZQrTgvnxkr/gDN/Zspvgq/
FVnAAeo7RUGGB0f+p1+jSk5OzC/VvA8XN1ifo6nL61TwBl/Y4hbrNghbr+CwphYU+wKsYzjNl84W
Zdy4NF6+G2Hds4a+SVTK32FUjKYzdMxQbkBUbFfK4PXwUlAMzjB+fd79qJcDM+6OudFSfwIdJiK3
JKq7FVx+MGJaBU4VKZfcDLsOSufJDWP01ktzDvlYeqzY2ijjIONZpFh/BTi4vY/gS2HaA0XnxWt1
FCIAGP42QKf1yieCTkI34Cl7j8TwAaD/OxVzfJj+l/ELY3ROWWrvGAoDgp87bPT300Ybtv/tmPfZ
OGrrXlARopmoeYagz4Tl+T9w4Q8sAh7H/vFTT+xhuZDaBxDaMW2IyGtZodkef9CbwMRsC8En2i3q
3dmdoG3Z5cFWwXVmacDGZmYlCdRxrGRLAcnxqpXqqS5Nn0EvJEjLxw0eCPBIo6SO1mTuYWi9U0Y2
ePdj/I/0VC57JR6iFgWITOQvEpK7L1J8ZEvL+rCFWpiaTO3mjSyC9RghxLGUEA1hqUQFGLIyLuJ4
HvAq1gigfaQHkBNN7v13iSUv1dfpVwK7i5cCiWa6Na5J5Vn5YZZP998S33sqlafwdHIvCv9vMbDX
/C7G2PrXfCOYNjLKOgSLMxC5uUe7pQ4oek1xFnDY8b89hJ9kei15Ov8mAbftbikkTw6YbE5WvS3I
d8mt5cpIPg8xj9oQbvYJI6wXnHMFCq5nxgYaFPcBYskd+1Fn1t78OwP7gxPaYFS68wcFrcMGpToC
hetNDJ/bvo0eD+4eIVob77c43w2bq9y3f2IQferS3wfsECM5r7TRY/AGfpzLaWh50EqnRuDozJbM
NPVevpzQZid3mnTjGGzEMyFabQ9Xszl13fjMsj6yl+Kjej8YhXmVjdox1n3A9xEPyHHpdwKhfWNh
EUr8K5YpQKTQ1XJACqMyPOa/nsYTqGAN7bHGXR4JvvO7GARRAavTt6db4+cch/mLHLSOs8UWLZ7e
X/M+gXj+HX8oIVdBawJUMfoMHkNJNDMa5eUj6QAqKG6x8WMYwwVYZnFRAHebvEOY5bFmv6BSi5+m
zm4IF1E91QX+k5e7M9BFmsCydsYhqv/FLepTWTC34uNZ2MB/VMSqX0dmrM8mYaACIbfqe2uF6CcL
eKsrv9XRfsRqZzHtVQ+jXxLvA3pUqF9CEWmYLyS0yHVlLe22H8Yz40aVDmgfVsMycJ7IYnxzra0c
rnXPYuatB4J8EP/EGrmoQLX+i9haZVckyfJIPvmfkIV9h8TVVKQ+k3MJ1dFzh1JxZEtzyrTIg1S5
eGEcX+7Pvjg6l6zHUkViq4Twd0IwregCvTCjxhwygnJPSxtTFSx1roIGi2o8yoPL19AN7KQkygrp
C31ek338gOMsDIB06TyoKvPkq4k3S4YuKHj01p73m1mgYbqam3snpR8VLzxEkD+6iGMjC3Jnh0lO
QLRPsFq5DoTZuvriMSFHw3Q2DR68r0H/tiVuvbwAnQIQkiLdICgVOtovfSJeDUQ3nskPc2OyQS/v
+MoD2dCWEBClWOwZuVRJrNiOJuFP/89YRvQnhlF63C257/0b/dU9t80y4MK0nDa1nIUwElE9uySd
2sC51GluyXKBlakZfpX9E4Y3Q2LmB+329GIJymYqAKmDNXVcLTYgH7dSEfslT81r1LRL42rkYdPI
mrnjFr3ynRAwCyJ0w7y6JFXjpW4lFCeb9zq0VT0GZWXuUK0M8/3I3MoMVgChNfsFS3kc3tnUaKbo
aq5RE/8k+hcxcmBmqQi/BrxZQAg9SAOMLapDH+V6Il+gFnViTldL6n+bOa5p99EU0AyBeZbLqmT8
DrJXj/3aUGhDvlOpvrRjxpDV+89XD3CU5XBf+WGomy8STCRYZ6Nto3OFIqb/jJvQUWbnpx8fhJGm
9xMst0ZOFi8wJRfhOS1zXPwxuFpNAnWQXJkegGX/o8uhoqLGbTkJt6kVoCnVsQGjwFzLRccny3qI
kSDVrBDWkcsHh8ZOzzdRkWTrs338NzQ2oLLOCs/QZ2SasvomerTY/zQGyODAL2dowW1Cn5l0AiiN
3mU7knxlVrHPJuCViegPennWAILfnyo/Z+bbK7pztEZ0s8GERu5lb5UWH+kr+RHvWEPpKtuF9aG4
XIcWAjJ+pUgkmD2xAgs+fMIK6jq4Zw6xKT6C/rsATLrENu52qP2WW4SY+RA4vXlMtSBDXt3L5HSu
mttBQhexALW4kawDFWLX2dB2KVoyx7Sm/VtUjq6avGD2tSt1FhtMpdVRhjtyze1xheusQUhu8J9R
I1my+J4zuh7tbOHz/2TSzeRixApnKI+YowgUGrtbVyV7fszDVLfKNn2omL2q+wSnU46ywx9AX/Ei
tQl0y4ufcyhsicf0H3PfQ2vZ5DHCo8L9cgkIkUi2sgLsL8Iw/aCnjCjp3zkYH5RFkZGtnVL5kOVf
voe2TXMLXN50GvnybyA0awudGn27ElwDZYn9wtzkHapVjCEKO+5y6S+Nz3BSXwBF5YB9H3n9MLAi
+ddcZXHD7Bi9M2MMqRaRczHeFvr4+fffFB1rIOLnIzbQAVB1McVIW3n3SU2ULxZJu3QQXSsUhyCz
OyqhUB44e5ZhXE6Mp7pm0Ij9NUW7jQgR7d6POjV1Wj/stx5AtWB6bXrvJPaG0eHPIXkfeDwevjc3
YYKgg8/k298LsESjQL3ExXfeKe/5a9KLOrsGX8Ygiwxr0gAH9cTTdmQ1k6jmx4eQTeKboTbsDpVL
lxLwh80fkWV7t2D9gidyIxYVsw68lZtj5bzCFV4IOPoWyHu6YE7aL7OF6XCIAU3BHB8bQA9UgVjH
6YifsJiL3vOwcFJE9RU5Y08IvtDxKgkTdCnYET3Ffoxy2RwBeCXPWbHowYUinalArMqI05fvr4md
tBXQN4I/skP8/GCcoJ+EEetOF3nTEUqnACCUgVtFHijDhq+pW/dwRFs6iFb/x0W/hDMZNkpVIT2x
bb0SaXYkt6BpuVxLjjreds/UNormJe6pNvxjANBnxEHbns4Pvlen7eZ2oKuHl1VV8y1c2i21kb/V
/vVM6b8m086EQ8A/OYFqdnVqm48c098uco7JNbusr3oED4LwDTE+1SxifmIY9zutg8F0+oEJXabM
hdGK6toKxXFbm6lAxMy5LmdQfJifMkfb8NRzX641DYI9PFOSpe5xP1fniJ/GQqHHbOZo1hhEcJAV
1GO/1eBhZtxp0zGqcaCj8m+Edkjz6TLkhZMXc/2lBRw24qqoCDUwEyewHRlUfCu6z+S+mYP/4lHR
drWYSyWgtQEwKVlU9lCtUyOdVaQYbCOW9TCTZBDVGdozrEDLUF/V+hOtbVaxnhpHnOdMt2jQ9V0O
yb6grsrAP+NI/eW7gVoSKS1C0nu9SGWESt/ENRo77JPYuFuCbOEpqEXsHiMUbxSVohGbqZUd34V4
Y0ycQVsSkx8bGniBK4tuoitVhL6BLffJIQPSDbI9Jaz7/HWsxaLw43jy9HxrO77Iz0CNR7bj74tb
1D8OeaggqOcRFWI5qY9RDUuuwv9E+7Gn3GExiVJbMiTKZXKW59fTgGocf5Q0pFZ1ZzNxKBW7V/fL
ETAY6nrxGO8Uh+n07TP91nCFLJjrRJLs4us2QrypskMq/3xVjMejtnHah9YGj1bwjJKLfJXktv5X
VBH0agt/Hxg/6RYkL5oRQAUrFX0iiX0//5FUOrTKuGUgczIeC2J1AY/5dzD/AbRpYIltUf0lAu0V
U7FqBSjhw3hxNq7qrT5mUiKKlTs/iBBAt+1xMDY5XA9Gfp7O7VF5Pz3YkAKEvpVUwsKTrAIom6wS
nxVkJQXAL3YcAKBD8neodlBULuK2s5ls472iW5g4FvMoAiyJvOJ0o4KQs2aFkFLa17T5J32CR/N2
W6dyjliFQNHDGTSTQHqy+vksXYkwsCnocLtl44EmuElBE6NT3ps9MuWKx8miR4k0qz585MtJoEVU
ZLZHAbGb60wfDvMdnCT8UeFcNy1GZ6wjZmyBW1m+lHFHAJhZHSXKwdKP8d+vmKd7CmtfD631kpaa
sTpdJfTgtRoZYV+oI8jh9ZOrKACD2IeOPOchgWKK/9qwxM797v8oFHPNzEzkYugYerMD+xIhRrJr
zY7hJyriIPBQLF6nkYCf8hWj7gMQ7g414pyE/96MX3cWjIQbs+LfmYo4gmghBbb/Nop6x04FX8TK
x7tIovAotkljAMNogIg1J/Y2C9yg3waYvuXY/+oVpc6w3Ts03rbTUaR2T2TlSXnBf/Bwr4xwTjcZ
K7PqakuAzFfXjOAHU4nYKfEjo0ErN+tciUFZbsXC4tKmDVtD+CiZZsVhAMZ5AF7ATArAgeLdHRrq
h4uZVKfWtrgAPIM2y1QKNYjWiXE3i7tZy6QQBKePBAfQybZkLgt/RNuSkluNKWiGLCPnxUW/IvXW
HdmYiaIYaQefC8cXuAoyZKNveZrIadVkyhXGpFIHiZZGI0z3GDOZcL9/wzIuofbhM8H988F+J7Un
AulMJuFH6CF2wco18xCqvhMzMCJtXZF0/fNJYVLdpJ6vefP1xu4j+HAsFZxgT+iIapbqVEImF9vZ
nQJzUKEdj40pQtFqbZyoa3hUPMPpU6iANopNQDM3ATbYU4YNIrnNU5f0BGUuOgEl1XE11Vsfw65u
g3BBeg1+IQ93Nt7+WozSWNkZWTtLXG4Ppcy1iD+p/2nykfI+YjoZITHGbZrktgf5TRzvDVQPZkXy
Vnw3iWc2tXP8PJT2STkfK8FDuinzc/TT5FKPtzWmm0ou4A/usIWDQ3PlQ2WxnXwCX7ajmmW1UyaQ
UTQw2PllK9E0zXhO3zhXlRPEH34KHjYA377wsDOagTN36v2L98aRMARsrfCyX5ZDwp+jzJiatBY5
5qmsSjf4RnW47vIPIamCOSHqeV0e/Up9Q73p4o5befwjnecGBIS6sLv3RsvCRzBkqbrAIHKIXXMg
sJNkGmquLEa54tUTvcQ+E6fzW7dLw65YxrDgdfgKhgDCl7cNgBGJB/NDLUB0WryMnvKzy8iMnQqP
Y1ljJW8ehbINV3Li59HXw7CYmPZj0bWcIXwjNuMYFtWg3JcwJPB7PirV57lsfCSiDPTBoLPb3YAc
3hlKt1UZw5eUeY3gZ4c8gcMkXAddERRdQvBpVnbrPb4qmDRk43edF4j/SrOBPFmFiJmB8WrxEQZI
7TnsDYlWFUhnOjaK5GXjStSPxYAbMyr2Rz6/j7cZi8UzDYUrMLSadXYHbORHVFDRxYlFjcIWh3s6
LmetVfnVOVp4MV7oogMeUA48KnT+tlJcQWebsFAOHHpjJKx/EKG3rIC4ivJeBaSzvAmQAV8zbTtl
1xpaXpTRSTC6T/C0T4523CMB0Vx2AAnelGq0xBOb2gVInlPFPmuPMwoQ8rLjhtMiM/+/69ZnaMOk
HTw3sdDQpulcn77Rp8s1eMGwX2X5maFMIJA0LLRNuVqhZ2oddbPuS1K7k7sZ+WfNWSmeVWn/LE5R
VDRNAP4U6M/BruogHDJgIJsijqPUde27UaIU0qUsrLfH2NyiKJ53OyLbWfLlbImU245o8Z5R+jUU
+rp+eqhENCO5wgBc4WVgs3AYmcCKv4KHgtDiFpKDqB0rBw7um4diue8Nb3+s8VV38uYLbRgUEag4
47wJzdPM9McGzPDIutmve0x1KcUcaCzrlp/ZGEo/9vYYV498BpjkRWVJYMk5eGLMtdGTvbtJC6rL
M0SHp5hTZLBDQGye118JIYlmOH3npnhEqxkv7dH/otaO9D5lq2jznz9WFPzJqVACnyZLJwMj25Ip
TJWYUFJgpi8tUOM+6FINayridVh5lMdcKG18t4tGWyYS6/ONjYmTbb8gm7U1fgBx4OxEBpGppJP8
n4OkTtrHQuDfX0GJz68IPmZ5N9peNHMk+0YCyMlGut4TP9V6AItJfTyDQsBDNOzQtgYkhGMmCsWD
LIavTbzGnjfV8eHuZdG8bCDXM/j7ok76Eg1bNTzbJJIHkax7mDi8Yjl7WUeE+1ncFRSZnVmmVIxi
NeHNrnkbbMMLVTgV0uZDgV5cFZWgPjSEcKLl4NE1JmDJvShHQnMAp3mG80jz2nbcV9aeFxMNqW3J
NjjSnEqwEnmtChyOvNfuUC02CK+VOr7Fm8sdxBHphE+mdAihWyF0GF7VLoDNpJIFvZ0RRZtW7MRl
RTCKjAbSNqWAtZlAnnUHOHd4xkBQDmiST/texHtjT0KxZYeXCCkkMxMNP7x1x1VWvhsKNIeFzPWG
Kt04fIE7kMk/d0dQI3m0qAKeOVsqgRpMzdb/pZiuCZxyq7isCGU5C1L6jTJQMrhHkbgvMGlahjqa
q2euMYw985LVQHpbe7MpAhNVW4r2GaQszMpywEdTANDe3Bel3hxNp8b9ZgW0pl9h1Dsf3+aP865i
oIL7Qt+uHFpsMfehw5cYVqPj6iKaW8T5nY3Z4xqf5MoUzwo4/o3kAMjywNdcurunW7dqSGOA4iH5
5pYtREHI+tm/NqRoGCDgw/VsQp3tahWcpcmqsuezHB5xskEXgdTwIh6hSBhkWAORT00yPD9OGUzz
1GVpDTQDna+m4lpN2Z+aKRCgQYaUy8Hr2zE76r/tceIpg2C+WXGtSKJj0lUze2BjXLEGegC3EXuD
V3+2vlLSB/k8iXn0cgvUvDqOmw0XA/WNrq9KGt3wVfgM7B7Vb7YvK+UT+uoP+tTfaKkPrmfxNo4i
t5BYmO/luH2kDX6uZOrwuepQPkPlqm7maTu5MK1hv/fwmTpRT5oenLqjuk+oJnfeLwgkAtyG7Ic+
YVGQZg5MBD5oP0VDMib3dPH0rpQ8xA1DaAgOtypY+WG1Oe8j/Hxe/H06dOtDbTy3OifoYZDcRRe4
g865PZh7FF4XA+9UAriRkxfsTI1fKgYKLJEUEQhev3VAQmnPrmKHQU2IciUR4f3SkBSjhBUc7DAW
I7myKyi/+OdjfN4apl850uopap0RPeIIlUvXydliuuIQkZJ5SRe6KaMcqzWlA0d7uWJVDNTAFCEh
txvOtV0jp/+3R0dwzi31hYqBOjiUdZyX8BKmOpnMfXFn+raV1KuLfMMCFsTfSviJoEjmWmpFnsyD
6dTCOCYNTCBvlqm6eQZlJdjYP4/4FbOvwZR14UdDMKTGCJoVDkWcXhLCkNTb5IOoy+QjLAmwPFdH
1hNIS1WdydbdjDQZBz+dFsKqOC/P4xsYv9gmc92bf2NvlNSlCTliBPSx7yM8aXMcbJ36lwxjsekS
hVC7W0YWx8/Beq+nf/9hxATOT2oKdPiTQOOk8LPfLOo0iHIehUQi+GHNkTDApYYc3/iqGygfhaA5
P80Ti23N1GtfrIsWccH0VPGE+1FXZJoQl/FfI5umE3PHj15vL+rFuJcPENKWUkHxsVvs3LyXssvi
0ubIjYghmPZHbrEClBZ+mN/kAMF1auZBEtWBo3fzfOilN6UP5a5BAFO6ouuoIKCzmsRYO9SVYoMo
7w4SLj+sLSQbdrvQbAshK2zHd6oGACRify2jHNkoeuYvnxc3MjrMDo6v2enBeY8AdmdJOtytGuYd
x9JsShyJbeWWuqUR8HLILn74ypII1ShZkJX1KAm9exNc/9e9B5gBbTBFF21xcptOHMNsgUuclk1Y
PFTRibDoY1nk8V7iq7QCYcZFfR3BUms9pAgl67GgxftsTO7M8+4fBLOVjgeGumemkRUd+5qSgeFB
E1hCdg2B2O2P/CFVH7o+30RRNkeDwkgGbLCz1ijONt8rJQJLLZdX3OP2jp5Aa/JnL7UlBhEZDYZs
HKx+2nftO9k55rEU0+Iz2Gq4TnRE6QMu5T08X9gEmGLUIudbw9z9Td/Ym8fkt+MgrSKanuoogM3o
lT82a1POS2Kktec1CZVgRRmZMSqjxm+SSnjnSHCy7UibBb2L6+n9n07NzLMPG3q2nWSYV9nqAdFr
uaa/KF49aVBfMHhGlHb4VcrF+/IfTlyedvVKrnLW0XmPjpujQ2qUB+mz76vSaFkx11fjJIi7wypW
FeijeFlvM/3NsbrhAx4foKsmsuu3EHB4ZrJN9dZWu71dlKWQ1sc1ID7HJuD0G3dMZlvj/vE+ZRRb
8/BJMbg/zcmLEFRWUWsulathfP6qxjb4JxOAl6Ohi9aWVBzkbLGmB2Tablc5MkwcSrrQEjTbyyuS
bc/pWdXoEpSTVWxVif17JAZ91kTTR8GlM7E2Yy5JSUzQqvydxqyLJcRhSrcgyIyzPdckomqZ4G7N
ILKEIQWgjHUs3LNKYKzlWMoVnWvZoSHWToLB4Ga2hGc5N11LOLzmHe8frh80nQqyAIZjSSI+5NG6
qTrkRLGSRbA74nvPQQcVS8jCMSvubnA1ghWRELyM0a4T5brWoaWBcEYPQ/FGxf74yo0WxyB+c8aZ
MDvxeMuOpJyLm6Q1HHZ1N8sz9u76XthRZQYxbvTOOf3Q/ZyYkPgxne/swrYqF7dzKKAiuMdzCanm
dQ5hYBxkT0CoLiR1cUvntDtu8/pEKdj9sbYCHMBrk7N/Z/R0glRf5bXSTcZ1oDixUrE6hhOjZeh6
71ukXNUWIupH00q61lwc+aX62YEy7fgBnimprQEVmTv4hV68rtZaEzvPZJsHr/EP3SpR89rmxgq8
9eo9G2B3a/twAH2caitkoQgSx9lPHW5YeU1RNeBU/T6NWrR02JjaGL/1sN0IS5a1/nYKlFuIQrpe
vcbvDsr+IKNuRNVZwlTP2EX7jI8XR7h6yrdnXe00AIWE059e3zxAX3u57Y0NTowMmViWg1dVNhgP
FNFPL+qKetI/XBdtXXxXmHkNvaVEh+BOhdBmUGI2dCgE5MRpJhJAQkm3ED5uuYtZbzhON+R++ZvH
SDmOamcxg8s7Z8dzu3Fs9N4WUtCtzxt81uzO85NjOpTXLtirn16zMpPjKuPHmNOTmW1j2TfpsnAg
VsAIQgEamUmwPZNVk0V1ZsG8lMg2lR4jXUuCE7u1Yb483PNowpUVHUvcT+cgj0e6hVCUjzpXooqQ
XlGdQfc8K5yyUJWvQGCzRlF8pD7us+dB5iYGduy3k0EsnJSuWEZdwI7h8xWi0EhwTdN0Vf5BJkoF
zRTXT9PbQJYOABtzIPzI7BvF/sk8llrL7TPSDRheX9Jz9qthFBd2MEirNwNGHkuX9Fagi2clH74s
BCpJLS4wbjnk1nOIsLuiDbi4nG8uljhjoSpRG8QUkmmp5lu6hkxawGxKuxpUVmtzL1EWMJ9Rz7BB
ZV2q/w1NgTj7vZE9vNGmNPX/Fh3436ftGSaKOTQa+pKzk1kGg2kgnTqlocPO9XhCLPGpN9l2zdkH
ZKyMYDsh7vyYFXb/MYpDDw855AMqp+FXL0CO/GK9PAkgDSSTzdu3/ARgNqgK4dQKVxgVrHWZtoA6
+IOdozAEcCEI1wDjJ8D5vQL5m6BYqKvG89kRoA7uJbH5UT5WBKvtqi4tY8ZZ5f1u7kzYSxvEh74c
b8LP8IQvNE2BO5W8jdAv90FMEbr//8FEvgaQW25uMGmwwZ2YPbHfbQLhkxNcB9tus9g/pxBR53rv
9ReGRTrjv8/2tiWrafhuJzrF/8DclcP0k1hh04v/qlejwpZ1KflrR/UuFbyjw14c9CK9PEBr0wWU
++St8jA/ll8ntHyMtsIbk+kiwoH64fTDV4ev/Gxwx+Rr9TUZIcRhVMtzuB8OeuEbEj32dWr+03IZ
rrmpKLSdJdvvun0/9I462utw9jhEp9GNrKdCOjhl/GPdyeisJ/M33HZUOqgf33yGS4nPL6nL/7ci
MbSy9lzCSQsSNztJbJnnCjb83b2Vu1jyMfatSPA/7SEAXfzgjX8LC9po2buAIR/k10olIwcnI8MQ
FL3yi+AGDcMqZapmzo6f3v1bMKK0jU8dSDc4AK9sh3ffqBzFcx3uzYfk+b2tAYJZvFfMJAWvg9Zf
9Ns/We2d1PvO75DSWlDrFJcJy8Vp28eM+kKtZqI0UTyYkahSF5LWJZtR2TD2HGPsmTm6qMbUTNpq
ARhmSOm1RF+mafg8bXl+6WUGi9BlYY025ILW1UZdJdlcLQ9Y7eTE1FsAUpkXOTcz5zThKmxp3gwB
4f2LtzaVD3QLHPhZQWWDLfYBzaCdxjt/pSgOOeK8crF/lPw2EwELIHAlFJKWk9u0439FT5t38w5i
L+cqHPmr97LkK97nARDAQSO4zpMlKipanwzl66O8FRcBADBJNkzMZ3zIdGrbS52FKXWKLyeP/0q8
PS1t3cYwwbt0dX5WMDfhOBXVGF20a3ncCfZKsh+1DNmCPSUUO09Wwbcpjf63tSQo1LDeUoTiSudT
2zr+XEaSCmBu0GQwjzRq5dHqOa74aH8x99S5DMUh4hVeCOePChNyzRQ5hVyaJ5LUaldB6W69uuHE
ib5ctyPcpr/FJZidGr7TsYivfaBOrFc6GU0qseE0+xoBh7126st/K117uYU8jRtI7VyeRoxuPDiy
b2+JTmZeZfBIX0ZkGnzbFIr3/mysBwbeiA4bVaYoqTGYJnwC3N3svDOH6J372LU2u4CrZWmow+Oo
sFSaWTtFM7ozgt+jVKJFo1WD3NC2GRj9n+gXs8eMiS3RT9nhvqHy+9si149naVhYAVcDhtsTqXgl
uN4vvM5yIZ+suRrPKW+sAbNysAMLadRbSdIoHc4SJCWEljLwmHVq3I9MW1HbRRvtOKNxQsPoVMmh
DJ7jnqRi5iza62sGX6OYzvhZMPGvPaVyLpbNs0qz50zMxKaDGrYHDZU91lx5qLdl0O32dg0qIGmL
VlmQ1ndMEUfXr0q3sf4BNCgB4BVmTU0RfiiOtJ9b7Va7IFnu3en/ZbfJOzww0/iATnDHO4HFtD5m
IMvE7HEa/UMylJLeZXkv0osFpoVVTfDi7HINPI3KpXhVqjWyuATcsbcwsNR3m+t5tLEEzJvshyT5
hD87GbdAdVKVtE9BunKIpssKSrj2PJ7kCy9u498p2p5e6/ZGLwTP+FFkutoPUPE7vHX6GRfQJHyi
bk4qLO0j4zFmp1KB7VpeIAyNSN0YXR+zSQp4zmWfQGLrkh1TOj0yfnlttfxu4asywecqm8LfMfSX
a68lIN2JKSz6SfG070vB2t3dx2QRpoR46DyK8A27nVgOSdOGbQb68Bw7Nsqd0D1Nn5K1sEyKIaPO
tEKrcWfsFdqC7IgmjNhKLFqKfEnj5XUMNcllvM9gtbb9I8pyVKeX3uqu1h7QIQwoL/I6/zOy6tbH
Tac8KBxX9zoaBNu3E4tBQ/zdC3CyFkx8bWnsHoJ2dOkt9vegRRDqa30QsVjPwoLNR3wepE1jaw65
9RsW7OUEdzfZ7Jp7RA9Lrb4MaTZIQk+CDxL1YGOBLJcdyNVw9t59LxORzS2cqhkR9rd3gJZm+p/d
IcBnzuq2E3t7F2Q5K6Frz7wj57R5DibCYKyRAegduNWOUgfJfzd3++996+NKnMPdfK9BBRjZ6w7L
7L39oSV3k5zIuZMhThae3FP3u/oyy7OctdfaKxs8X+OHT14M+Dhw49MIcT/y5UPitHWjz3UREmj4
FGWo1dUCKTuROI/I2PDci6cqHO4Ec8fPD0G3ZAAnIAqoIGoxmC3RmK4QHpBm83zX6WZDPSKeBgSJ
ftjhTKtvXS+iz771NMt7uTLpBkcHodOuyi4sMnNxcOorV/yZkf+ObaP+7Z0WqPMpjn/0ROzENeX2
MWjbxAdesDnr963sfmKOSG8gGQInktzRELTKRyuiy05WTq5OgkuMsGj0ynPxp6ASMRiF07CxGwfc
F1kq+uezbvyIWnsP/HZ4ZVIwY8BypjIaVc+UoJ5pevE6Cwxrii0CbOs4tQhlCF/TutA64pOKK417
Ker1l4VkopvNyxN/cqkWmVAGMBWYIvfnqc7RSxNit3YL+B0f12hIjz+vG0OgXtRAyFARdjvXXCWm
JWM2FB2ggDQSFmBOTNa/Amht1vl/vHOjMxwDsAslZVo+RHkggCnmtY3uKpmeFruwLZqPNSjkrIzA
4sAvBKLnsu10z0plAqw5Q2FwUgPmHE8OkT30F1/gtpqZa3fr2Fkvg+XuJEreJLBdmxEZdDBzjNO7
VY2bucKTnzvlWUUOORQZfqi4YEEjAOIfas/BiyUz6/Mel0pmm6+J7BSRUZXVUWc+E80q+16r4l3Z
fTKO0RespOPFoC+2355bGCM5W2CnJkMHrQ5lEWredrHRcOcxs4CXNDtxAbrYFb5agV0cEVrvhpcY
o/M974GY/mnD1fH7CjEk00st89KEYfv7Fn4bge/hkCT8UZt74T0DocnFiGnyL4s/bcqLLHiuSvIj
MZDtC8nNx+9qpRjB00GGzlWLJaBweo+3z3rfuhyLELwBH6TAB4j90F5dV9l3NKbJaW6TWT8UTYfp
tf87LBJL/R1vU29Fg5Ltspww2RvHsIjGMXoRGtCJLe0HkmynTxboknUiVxYmZpLnz0RagqFZ/kXx
yYow/eNZCCBg31JEElUX6lmGx5XmYrcQqD9oYwDge1XCwkwqOiCWm2CE8OKs8lK3Q2SAbqJwhLW+
eBC7LcCrvtfDFJFkH7IM2GsLNTB3gPF8j/n7nwD9eTQ8jvk8MfQNEjLocZLwvFZC2SivppnKa4EX
h3Wi71X529JqOvuz0sOggnFilD3MYLxzVPRj2s2hRs4ooCDYpeDVEiiL1ZjDLuvr7QKpl0l2wENQ
xxMqmuKS6v7144p4U1BWbTsf5FFpSJp1xDRzH99icXlECGR0SyqcEc69/FUM2bjfspQI7+lF2YDL
Wiot/4YXrKcSuulDlCgHZ04/CStzUemauq0iCh3/R6gcp6fVKWh5Z7JePYIXPv+FGxUNoP1b27sd
rYbLrlgF7WjDAFSUWFi8J6Gh6ItzEi19Oq42mrkfqF9y/TYs8itew7Hb4QrlMJBXcXu7KGKNluAb
F38EqRhdV1pbA/18lckhmoPr3NuMtCaz040uuWDNUdjnk6Sk0BKpNUB+VvgFwZVOHJ79eKr6U29F
fsWAh1HyV8hg6vDUd4QFdv8OoJWB2sUuy/u5/qDnyU57xUSfZrkU3TFWta3IjjLt7uoqAHGBAzTx
C9HqqA2Hvhjj1/0oBXdFkH+cyouA5pI0YMMhlvkdbV7JFcKl+EyjHE1LL8q066Eb+4gDtAoL+YC7
6IRHo97V9aOBmW5+BJi+G1g1FjFODOWDHi0CzBPxi7V0hSb3u4/+nWqeG2zodxjCHi5GNsIIMlyV
Sv5RjIfvP5hHODryGQ+Y5+g8GFUTerHpxwa2az/iJeAvpFssbl/0AaypcrAa74XygpHWRtGCOtq7
L7Dnk5qXGx7wmnhaqLKljSDFy4+ZO0pVR9a+3b9wN6eZwymsAwJoRrfI+ijxAuc9j5sbAEuHWy/F
pK1hGxt/GSKfXl874sHMkDIj9+XhEMNRRxt0ZYJFSLKqA9YhPWBNGLcmzLjW2c0HE71YyOnjmkd2
KEE16ln9ekTKjVX2E91kAiG+CFDmamLq5bcmzOX44EUxlISnGIXKWfONSUTLa1zuP3OyyfVi+pcr
Qv9jBpcZJqUuATCeKv5QKaZlz7CpvcEImIFeI8P5tT41ij3G98nKybDoKD2OA6qB2V06Izd3/6K+
hfQMhV0D100BGHGMpWN091chZF6eb+BoBlNSox8hSaf/LKMFYMdZe3jmvR5WNwkGxHaCVHrGp9bo
91SFfK86k84MRgMn0q0YHUaIyx19VOE41pK96HNna50w+NnOMKokLE2vNMFUDtA3nP5LnqgnKbTz
OPwzF9YCOfrebQqSmhX8QX4YoUSNdxxMmLnqxDNihxK4+wBCgPZaOxyZ93TDT58Z2dpERe6yJSot
bPcYVW7zjnkHzA3bE2mxw0zxQsbzXTNaRj6YiBl5sW7TpYO7YVlgPEFBkldw9WjD3x6RMp3M0jky
ZnqOSJ2N/25bUl5yRl9iZhIl+Y3vx2hk+L81jlVKgXtls1G8JPfClf86HxVjhYrk46CjXSl+t8st
76waHA4BqxMhO/BLdtkAx/+whNCSRCcgE+U+4Bzy93Eg3YwrXmXEkMaSyKtYpuRqWDoXnDNnNihh
0EzRZqYhFmMRlNKjSU139lfBwrRor/24CErArSLYaQMcWRZAV2hqgRQ8ToROey6ORcdW371SS+zB
Oz+w392YuoytfXGoxQ8vMFPriIdyv7avyeDnrzUByF97hDk0yhOtl++PHLbOs5WdBb/s86mLW9Og
CDVoVCasMoDHnEldG/yB+i5UQnOs+XcbsuJtvVEWEGgojes2Ewt6slwSis3KDTdPqj6wyanEmpjb
jzsp8s+yBSP+fskSEyNdF5gMHXRrvkRTPRHvIAR92PPOwASoZ2QW5JT+Ovy/poKUp1XWRVSGq2kR
5o325C6QWtD3zpQ1vRTsSJZknB4+DvgpxM0uZUpajxU2hT6IaSRoDK1wvbmiIz4R4n56EJsulPCk
8Fr3eMtoW7EpiyOqW22T1bmnNl0iN0LIbc4YXyI8T2fPCaf6On6YwNBspeprEO7fhY/tIJwVB5mS
Jws0AhjwpDKBIW4FW54oIi9j92Sze0z02SMHBYJZlhgiZq4DMZaw7rYWPUU92n0+eJkjeS3cXAIV
j7hLcY5UWZ/6lcaq1Ec4NH5VULoMMwjrRNegrXP8oCc1mD5UE2dfMTzx/ypBs6wbwjN3pHvuda8B
foUK2LWG+WiDFBv1/n+8V3G9GQbMI07GnOZv7UA/0JzkUnkIHYfNlNjoxEKApikjlgAWWTExwNzC
oM/dz6o1HNHobXuTxT6tbAeAyuNd52s+M/OC1tl2wnP50i0T7BAQHjezAjy7sFROaSzTTlrH024K
cLIkTH9CgwbjciU7n5RLPim1vvTzEguGipclvNykh/wmQaYCollSLhSDR2fj7A84sNt/UyGltWtf
xtnWL/2kxQqtwhdructaMdG8V94kTIot3DHB+RuaChsibbDPR/Ke2UJsgcDBKoFM8pymoJO93f3r
qYqEv/Xs7u41Va22PCsXH4IrFcA0J6WQIbxVygnhlTvWNHxOrTww71aJuD1iVr/dFMVHwsdrw+N0
LETeMsGmWyRUtWkaW9WF7I/403jEgfYh+eiVLhSZPAm+IvK4eBNh6GdJQmLGoLKIC26CtUfjqbQ5
5x8w7XmaK6I6DQsbyjv5sB9t4lSFeDhSXFMBEQm85UzV2G8vBrJYH+Eu81pfcGCbNGHjxXEdx3x5
G2usyDcSiG7lCoJycoLU4BndoeU/WrdTnUCyOt8gRFs+2LrOb9+35t37ChjwldToSP4n9lSA+oyg
lv5wWS2QgTid0pHSsROTiYQZ8AtzRd4e8+hjNi6J5Mj40EgY7Fnhaoehs9xpA0Wek5ASVpdJ9mAu
JfZ1SJNU4ZzuWssPeev6PO9XaPeLQxmrcrYzBAHZkNhZeLflGoocOTLUFH90y+y+9o9dLT5bU0oO
oXV9BIoGBI6WpdA5+1geKuxeuC7TCYU0LHrpSAPnenBU5I73MF8QkMjNczlUOSd2GW1oB+KZa3wg
/zilbC2g3qJi95r5GnVBTMV9SMRPdkgCac1gy9o1Ny8n0bWNcjVGbS4I6RiuNkAOSDc2TJLnRIhi
kFK+8fQCGsCH6d4nf0OM6bMnHQ1JyvewFEjzptqEWCWkzqXr263rfSHy7VNyRysUS3lSlvUcpky4
ADNaz4MQxXHKvO23jKvSkQdSz3ogUqf6dcHJryCfzJ0ujQFpWDNH02VNnpcU0g7uivFTRAhWNEzj
BDmviQ9o8RoDhn4611YXcwSaW0+Vcxf9d4W/dP8c6+Q90LpXTfkc1URNQBboVUwA+nLLmMSLOS9H
TQTnaSgsOXQWt8lSN2HSwUlSq4pRcP4jYYqZ1xUG/5xZcAX1ukYhGXrCw/zGj2OKuFoKfN/l0QjP
uFpEfaZVKlYw62Xi+puyIk7o4NNXgS1zKHr/DtuZJNNB1V7am5+DAHii10AwpwFEYeavy9WpcfbZ
ZrJmlnLBUPKMh3y91YCU/FM3Ywzd/uw1hDrBOsxFTsilYgnsFwzC+ifnh5wwIWvkDSjDd2fsWWJY
tc1GHStMzsWxoN/YsptuyNhjIwcgLAf3r+FuD31zZTSaBBWQtsPvTKRInZ5vXxIRS/zwnLOko5Qx
MUrkBc+AVtX0UwmzNH4M1jwXSYBQOdmIAmTxokDeQrCH4D9HzIK+DHNac1AEmxLJT4LE3/EIGfgR
0g/nWMrUm10uVhVRUgKn4sQ3KKhk7tP6R6+FJjFPAYL2C24gv1aMDbDmS02i7jSSR4XFkHLfhwPr
aPpGAP/ZKZ3LZh4rTBvTQnI/+nkwYaCSh3Dr/oZaD5J0NjqRBSnIkDanUgIuJh/xQGhupz/BOZ0o
P+sEosSANkz2y2ev941x7sF4mDnYXTF9j5fnjnGR05d2MriKd0SNjVPb19oM2zcebDzjzFKmLcY1
SJclcJ5l0tlN2PO1UjJQ+5rz8/DlcO3O7K8Cs9a1IJgtefgeO8UeQ+wA0ORYqhKMnG0JWtwH1HX0
KZqyPi/SeKlAXXet9JX1498N9fMBLjXC10nRQdHW5u+WxwCmF/S59b8cvU4M93WGhgtD75KU7uXj
B7DQ6tqk9+0xCcXiCR2pjUxdbsb0HJsDF31c8uwj+KMKU+Yc4cS/HW/AxPsVGKya/Od6042K2B0q
Lu3QTkhlJmqGsI/ooO4LPD0WHsyAQIHVOmsliTgvJdm+aZIlZqI1NzrcjKKK1OGwGibwM0BRcEmt
j+4HilTsrs8elKjWiDth6r95R1nfJ7Jbb0BJQx89NUQrndW2jWL20XfsN+OrkgnfcoGsarbiSiZ4
r8BT/iVuGx5pSbmomI1jf6KKzJumrB3TbGElrPpFLdxYNFq/jDRMm2kuZEAmKCMFR44OYTGX4OJ4
lMiYZvD1FwN96wg1qe7a+hoCurvGRkDualT26vkv9GalwLIgJ9bCm/wxy04036Uqhjzg1qKbFa3q
9W3fSjItpoI3Kid4NyG3r/+U4zKnfxdLns0aJBw7HCQB+4/30CCijapiy8R053ZqhlSUbdpHFsUr
Aw0g1oCCp2g48wzDgaleoY2mVtJUIJRoyXdZ29pYewPkvvY8Zif2DXbqeEIm5hiDQhcFLpZwgH4o
tkAIRDIo+xqi5TfxHhzlTqspy36FD/TX6Vn2oMDV6l7v/jbld514rSkrHFkIRzr/i2oetjJ/Lnx5
Ne5KTdljKQNdrOoNlzdEUx1DB3+LeEtSCTq7WRDnHT3Lrx0sd1XvWD03YzGpfOtC4VRbJYK5zYNH
zFKv+hZlF0ENFnZcKEwpotO7ZVHM2QkYwNouot6W8F+30yfNlocfjRTy8r7KtC4cKVhfa6C64Tp3
8l9QbdvvHP7gZHm8xJ4+EWyg0Zg4OI7BKe9KwwYsAg8NYUmnPSsh7B6WWSg7mijHwLsmt0nBpVcL
wUQEFTy3noiZLJh263O/TIR7CFPJqSeC0efOJHWBp8ifAGGn3+Psqs2XNLjTIkq21Jxa4yMXV/h6
Czrahkrqd5HtuXniANrm7ulwA3+VRpA1Kz63/Y8Y5pjfw2EdhOKnLFoyoD/1/laPZ2nZvdVb7Z0H
p/z5QKmCQHXyKv/sI9t/ypfepi0pAhF9GqCMqYKBgQNdg+MCvVhDc3sevyb3MeJHsDAmygmJsToS
wh0TNIzT8fbc+t7im3/JU+vCgcHmSNsPjbzuD9a0TV3kCvKPFISZuMzN7wYTdIo+AeSbKQVTmtIm
OrN0Rr97CMgE+R55UO1d+sSJmx40Wea2sUAe8vkKdWrJ85njSyLP0XYtmtgwDRMFgfz1NzU7EgrB
+lTaFLhaFZUyomyLboTy8b947m8r1A7TdPMd6Y0z7pwyMRnqzRlShwrOmAsag7FZyz220yfuZY6r
+MFu+cVNbzQIWq7j9WT17zTSeU6fKNkJyvmKI0Ja6NeHVNvG3Sd4t0tfcKxod4ReRFkjCCIRNFq3
+Ujfq9a4zIlvSUxPIopYKIhTTc2/jeMWoEZND//L0v1TviVFIqoSFuk8/Cs5G+1jCzcuJMArck87
q+QFOQDcd1ersI9tZEz68lH+rz8hB4IQnO0dWZlrQmN8THyIs7BzSloqtLbGo3BuGVxo6DeB+On2
g09170aiBxZhK2I+vDSIpvHsqYywPWCvRYwlzb/+pYtLuUrzU8KpwhnGdT11zRSDUJVWFag+dCa5
y7ziFnjOTS8jGuc4DzHcPWNiXsY4dI9IkLspFIXP6rAQgaZGTsO+7/FswexW8kficIlO5wI5fbvS
fi2wRyXzRuxFPGIeI/27wa0XPMZ9HhgTGcHkbbed3DtJiu23uj4/WxkS04RmjJhi4nrTaI5XuRbs
n6Obo+FexS7UNA9vkBGLJW1lRgOf/Qh6zJ5H0vdv91HUPntlIy60wevfTu9dbmHUxVrFib5UNq+a
/jMlJ0GctKoC5swubWSpsihCkAsx5MFF9VLdg7/QYXM2DJAz90e/ZU0IZ7WIFJbIjF+NdMchaur4
15SWF03q2HbhcNSY9qjjcHagyhFYJXg1tnGu4hDq2NpQq9vKPZ3RAi5xChdI2Tvv4Q89tlXhBMCk
ivQVZ08WkDZ1x7MP/MQkqLVhyPc5bw+TSgwnngGM0u1YdA2sdUaF2V2Xlk8g2ir5xKMpqOJNJPdS
NT64/4mH09Zi+QZegwvlRDnL0OX+++JkCutuu1SK0a6E8aq7LE92GbMK4HBdGRgynfAPUcwdpNE1
wSNJO175vrsw4Vsqi1h9s8tzzOKnH6uVLR5hKP+2wY9YE96yv+7fGYrjyqenyxtvlNeFE2pixKq/
PqvPrqBqNA4cug2CzM/z1iVvqPm2WqyNbHlOrZyxKSHAILUfqQqhjL+xUr/WKq2EkJ7v3pBrUbBx
+QE+RNLn5EZF1fixM3fWipgnpDVGoWn4IJOYES8xQXPFbY+R8JYedYI5FN267VFS5pQ5tf4sTdRB
VvTl2uklA6Qxw42m2z+acX7X19iX12+wdHDIcNEDP3xPUGpwhkaCSYTyc4Rm4wngiHuE3fRtXEAu
XXdp2vGih1K/nVE0M7sgwO/JRbrguqTElwVFnCo9Mle0lS8ks9ZjUkzj182UDnbzkxvOir0GskvS
UQBVQodrsri7CG04GCmIsUZbQ3w+k1pesqFDI3GLDNreh8rfOi4vMMyjpssCKQhjpzS0+YXnXT+s
y1bfumwKoh5DcAFSVDgBB+EkMqGLMoAZLlxaR+YKscp3iJK/xJrhdluTQ28GXkO/sYAZOR+1A/f0
nnAdZ95KYsaUA6E/zWH+K/15IVelO0RBuJsYZylBfeX1nVkr4A7cdzhWT6jkumGJ/lray51xlxb+
63twpVD+3+8I9Zr6I62Iq2WJREfqorPrpKdnxF0sCzDZJFQEhj8tOSojFNTO1c681ijKm5uGL+WT
SGFVLhMaDnkfu/qGw0RHMLJbv+KDa1MJVS1/TZgEsU1dKnmHkIS1XK7gJV3IiCeHSSu5Hpapdmf7
sjrhIpgtpEqzaBr8VjWAq/B1Y56XW9VoyzZcmVjmYhu5B/nWmLhQPhibRKdMppAHjLVxQB/UCbOK
XYDOtJA00XmAfhiWhSu/k+p6NW6YYPiabNP33DO6J6FXm47GNu7RSkLO8Y0pGLsSCuqZLCgw6j+I
eV8FayxlzpoRBCzWKLG2Niwh6sGwXI1Ml2nhvF5d3Yf6s4f0gcTs2Nc9cnnmkZkYgLSnnaOt7Q0L
faz3YD3YWXrbAiMU7J7Wx79kyt44sKyGTGU+aHdHlh+7A/vC3IpuzDVMmeM5PlySMVkvbBwtdada
MtjqgYxKOBL6R0oP5GsrJ1E8Vuy6eLIske0WdDgtPHAQx5bo6UM/S2FDIo2BiOANfap5zPq8ncoo
2r7t521YRgR9lNOu9dLk0Tv/Ckwj/zy+7YGOuLJM6ik66F7uFt8FjYF3rY9eTU+RKeWvYPGkdQ0e
Skq9+eag3Fs2Swo2Q+FWostOnyhK4uRSBJE5haysiH1HzDg8Y0kfnjepAwAlFg5i3yMfVjF3/Wyq
O6/Cb8APc9/lg/V14r+5vkM7YQ3aUl2q1imZn5oG1HY9pJKJ/WlY3+3jrgmCe6tWQ/RW3ehf676m
zCKrxAWPxOfoHML+OQBUkWIU4wFDZRtLfakOAzu4LJhVcVcL2P3CtOvXzrqUoEWb9SsSNM/rlklo
MJTiXSh/FSMzZzzH2W703HzOWsR1PGuAi/ItbdNXOCN4P0g9KdtN9A4fZ7RKriVDcFts4k6BfN8M
FVfjgGmkCqcydVlpd/ykodX/11RlrRpwsHk4rMr2TfGJPrBH2z5y1vQdF/UZhOI69/C1BqjP1wfv
JBmie+U3AF4YOXApKrfXlP0zVv5SRpcmKTtFUMNQkuINLHHSuRzKQwVk1ZEbtj+e6jLVVDUsQB+K
0ThAFTRn3H27D/zOMYkeY0UPuIuzxzBgOXQOAa8VI0DgGmILEp84VxGb97gTXGY8bTxDNMoBftY4
TyYGxJu7gfFX04H/hM62u12aELlMqZ8SjArBch3nb7CCEqTrXD23UcjHDXY4c2MVvkA2Xuilba3i
QTA697wKAe3dKzuutR4TzOdSe4XvGXrwzVq2PN1KadRCmxI77lyk7uyDmtxrDgtG8xisF258r2jn
cG2/OaYy6i9KLQY0nlhUr33k3agPPuEt/rYWQ+9OiVXonMpHez+BHOwD58mVCFvujJkoeeusgsKR
Bs/P2s39wQQ8d2hwQ15/ajwRRxwyMTPmZMChRqscOqCQwOwyZi3OZ6WSCeg5f+ZT0ceP3eCjuCD8
Zj36oEKiOvlnGoX7p0AzS5NLh2SBQds9kYh7C5Up2VIOjIIe48Iq0mP2U1BoLkPEGaEcMzULQFyI
rcKReLD4PHNTJUNtwEKcJp7DpXH9+gxpyNVAgeCWV+uwwCzl/VgmWUmWVz4bKn0U18S3EaUFhsRn
a8jn2JIj4DOM/lXmMVL03isYuTHz8jj/t2nAADGaCh9QkqcYqfxt4V/UlplVGTbLN40a441vpTR9
yNp7r/okqJgPhF3qLS61JfJKQk1c6MMx7VUn7fmkuE7PYAibcUMAWJIeoPZU6ueOEqt+uXxtpgBz
GBUqADpDRjgkpm+kJ0+jFcOedHtpx/kT+JjDfzazLVYKJ8lBKEXiUQfJsMe3A8iloRCebOZygMeU
j/RlZRBJ2E10JW+Cx7mUVKaWUzHVq8/0WBOHqik8AaeEz34Y9zDEQatjqB/F64qzIznCnTZeL5s6
5BDrw8W0liT9kvtHoaeL98GO/vpM9NZsef9nzpBP0aJxv4gqrSispiykExObgIhuQ9nrkwH8Nqp5
p9d+IVvl1MfLvyflvyXf1MfdBZICTOEOoMWGnVLlXbLLFGrSFPEoGxHIx98Kg4V/L2IgtIvgzMRx
9trkaJmH+nmp4bQfKBCtW7lqFnFuhzCgN2le4uhPHBux85kDX/s7H0Z+45D5H+XLv9PedypjaREk
OqYI2EUo5QbAKg34SXeThMAgKGirDpiAehFVYSUe3Q0x1p4qJhQ1X3jhUimgtJxocg8n5IwpLqoS
+nGNl25FxZ1gZ4lENn7YowDEhdNrRLB+2d94hPcCamGIV7lqDHkb8FV33XFcdC0aSX63JpXrJ3qF
3U0IUuvQ0wC8WZtLFzATK4oYbhbNa2I3KC2YZgTVBJ/ID9EgySawuM1vK18Dfqz6JtOMPoRfU6Fh
PSwT8zIqkE6MS80AnCNhLmmGi2aonixU6O66sUIiXDhojZWIKqR44VoI1qYJooCgZhsJggwwjTfq
cBxnO2nScoWvXj9wBIYWJ4kClfKZQFLmHkswO0cLmqztwvGE9rMuJISXohoWH9Ukpfg8KNiIO404
cC4MFuxxFilcaZU+LOeDLFM8J9EwesmjwQV4xkWdYCqzwiopS96MUm+EUSWVSRMbT5xT32H6ujQ4
A4sGmyY+QRv3Jd1kk/H60l2DlknWRfqttSHguwEuH8x6trBFYg4c7fQJ6Poq7TxxIzFU7Y0Z4geD
ZoZc++ZjOc2zr9s3XEpCF+UHaN15gKeeIvtixcxhXsoMYObCLzFD0cHwA+KHTU4xpag+uDALohWU
bYj798BVZ2MezZF1/xhraaixOWzxRkyWAc+M2/WLk6qgMFruB04m7c7CwAq6bwaX+Wcj7MjDgCuJ
IoKAETebibgn1WiE7qNN17+dGFxy7ihoWooIl5M/u5CsU1Ap2ji0TsF46IfiWmHLl3AWyvqqGzeB
jPIg8GHReB73STC+p22g+746x6cYr5SsaCQMRVJOWE2yFP1qdMB8gQ+LwGV4FiR9bTszNfOTndx5
XFByx8KvRrFfIVJzllntncYrkaWUb+pPE8Be608Wm2NS7r4NHjGG2oa6Ku043nCXl/Dt1UrsQlJw
Tw8ecbidRyf+MkSEEo2PZkMKIqCh0mjaNlGrWFAhcKbkq0uD4GF6gSySwHB39/Gou3sjb3z3rshD
osElQBGgYtoOOpP0w7WzdPQGOsixmTlXGsc85VAh9lXE5D+1BHvhh1+EOZUQt2M3In1gBrdBCEJz
UVaQqPpLT2/trvC5yfEj/9OmNjLKoF/NwDLiIQxMjbAziXk5IqRFpLmKeWPUdDXjVGZCYmGMsZuY
MimZf2D7r5iHlHhc3t0r60B1y0AtyUWk+GWinvPh6OCyqxoGNQIJjx9qWGB0sY7MKpPrMUJa1KNt
d5Z5+qsRurIGFJv0H6d3LNI35Fd0vmFIZNqqKqEksUHB2UxJiNS+pgDHJ7xZnbPFwG75nH2Aw09P
VtSCsrgAnLhUCdO+wDF+yGKsE7nE0/tfVx+WQsciz9pfKxC35XcdfYgzAN8IHT2FUVgjEwxWCMdl
+auS1lx8buyKemAwjsjtFuozTzVpXEFKl8fuqrHMDGsoesQ9cJv4LBmJHcr2oEKK1G2wW8y8PakB
0WUKmDjQgTxHJ1ce+b0Fspmea2BhmfXpjWjW/iQ33yRIAeLzfIWxV4ZXU9E9wQYRPKokbsjrZX4N
qS3vLLcxgkIaMN0ygPenJk7I7GuYVQFv1T7TZUEH8MTCCGrxRQbsFSHLmb9o+9ch4jWyXaiR9Qxv
N63C0a9U1f8XiL7MWu5brmAcj/76xgv9Mo46WIEHBwIYtQ9T3Iw8mUb/Ra3K8erWcYeZMb5QCbjo
4uXxawlHulm2/W9VPitL9YB++WSjA9IWOv369oyoRpU0+0cDV60J+paqu2pQt+ZTfvTd2a5lf8n/
x5vvvHM5k6492/udrSxhjRv+cdsZZP90VOZfd3NjADkXujSE7I7Oo485w/lJcs2ve4Rr4WBz45JU
x7SpHwZNDr7YWtWrRmtpBUET3Jb1ydD8EdT+K5vsEfEKzHd65LJEd9lzP8XJxq08pGGG5L1QNjQ1
JHMildCdAJvfVf8zyZRWBZtSBMm+AxkpQOrCvZckpZD+2ON7T4ZDoYnT/shlxPjwepxKbhZdwe6n
sJzjRBdYy4UTWP4A0so2YVgljsSytrYbDn6U5HDe0q9Cfe2EPxXhLp0CU/p2t4mFfiqezRFcCUWL
drW5F0Z1OFpbUBafb2CxUeplX9VXIyM7zTJOfWV08QhziA0IkI/2VSfuywGIxsAlZwZJO0P1yCaJ
2MGDL8GTz7bdwRqJW7WihMnMXUpPA8ONeG9y4hn/lWq1NGcsnOZpvI7I7NjOi0xwTZw8n66kJa6y
eNBfhJD2ScFeDTFptFerW2in3/ENSnGSygTkIYTr+yzVZSqgeUyk66gAZpsJeDzraJpxbGas2ZR/
5exrinoAPdjsOvVllHIU31CJhgcbGJA4k1VbKAx+PEzZ1wtJTSW4yrTFGXC9QgUCs6Vo6GSVaPCx
xYgjoFSbhmJD5vkH31sdpFT/1LOBDS+5J7ECNh12OmslSUduKSptxpCg8oi9bQU4ZmDksSgZ5pb1
qDgCs3Rk20+4Kwj1uJnte0+NU5s39kitUyH/AIhMBG17SQoLxR1tQKCwh75lwJFFPFwsAfi0vXlJ
NeJpUuHF9Hb254eHOWzV6rU56ePxw67FTOFZ8SwK2lPAg+bKtLTQ8bWE3+apSZGlXYkpO4BFYSaK
4t0ZHgtCW8LGW9d1wWSmOr8xxTOxIIJgHKjf40LjmBMxNmWXV0TGux+ywftbZ5NTwMvG29x6qmTA
nIiSMS3K8lJT9HuJrcZtYyDv1f6fl5JvrL8FCKLJp5UIz825rhgSbWBg6NYVxQxw5rboEYi8rQR4
99Xn+WMheoH1lklIMWV9cMPp6ADsqX0pVAz3QT8lUIKVtC+14A3Lz3HXqWRzhRa1Y2M88H4v0WAP
MSfKZ3ZUlPfrQEyRvdQGPkevLNwZL/ttnYyPcZLYnvFf8pb0OkYki1O5o9ymHoCUJXQ4fFYOk6Vv
PWiyj/RLBFjHzRDyjXUrHdoNBjM51u19vKYhd7TjaDJOYJK6/EtzqbgdSQYDg3V9lCpPrHgDAAC/
nvarYavA3NjvY85XUJVxlPLdpv7YO2hBzYbQLbGKAMjVBd4R6h0zhTOU2BPqpZHh5uj7QCcQwtXx
lGTq4ZO9HPG+m4Zckl/VF2JALXd7m+qaxFPlAIbPknyS1PCurRaziENWeZvYjJQyFqLc4AAuukiD
v/rzyKCLn11wIoVKPrbDEOw8NdwNR/6yrCXZ6FTGSmkWrf+fcYxt7U2A9HbyCrnEm+n788N65kHG
wAYS7ko6BPOX915ocxCiGXXyBiNomnlZHWbC7ZbIegns/gaPr3rfKVBJ0cTKbKpi8aWq6FEYBpmQ
ZZUKJDUuKU+ZRZQVTc7Ww6ZPw4huUa3Wyi5gNV9RfewJ9P5lYK/sKZUwJLcxecfgfDv4QcFVSv68
SNuCtuqczi0mb/T6zHGEf7Z0MzGe4v7EwD2tg//i/sLSS0wtI+c1pVhcTvz8KrrObHfx+5yWXQ3V
t8gOdsrI9pDx8HOgW7IMFmwCFKTdYtzDwB01sX6UdtSycBPM634twfbxTR/XUf1zBB090gX8yeey
7yF1N/BdKB5HZS/82bcM6p2j9akyRkH6gi3s6uIRiW/FCtsFmlURF2hOT1fts8dyJVun33nuDVmc
w0LZkjiZPje7ylvQ8/Y+12MMF9Xqx3IKSjjyUCp7kb0H4eIaNTg72zlL0oqN5ly+ZsnrXtCRs5+K
UH7CJ5Alf0NmCxAT0Ouj4QLmp3GjfCK3q5/BB1AwdQwWl8kGHFrslmiFtTcV5LDMxUMOtGrdIdzH
IlXyJD9S3+NVE3h7EWVN9Q/vUs19PVvSMG4SSmvwjy+xOWwm6LbIQoE5p0JLkWhuNoOIdaw+mwWJ
v2OHdBVpppJ17BKVE8lOUSBCZyGmRbaYlPEJnsx4aAKmOHAN33XoVgHtu5mXCqYCWgLi6G8QT7fl
Ha//3DEAv/djMYt8vx0YF9+zWK6g1qLgGWQTuVoOlZpXokmF6laLjPqFG6TK89XUPwnT/0kFW8ON
bi1PIjyD17HYBSdBZSVDhOdvVhq9Shtw18seXAX1HfG9b8vasX0EbVEsL7mddDt0ATsnu46qnkYe
ZyBy1TO4TSGmVw4Ycqoulp7v6F0Vkkon5tOkzJzpijwiyvmNjQaRIxHacN03ar/h7EpThw8fSR9C
jeL782r9g/LjdjkxAWIBPKtOsYeGatqoXvumO2un4VZARsxp8u7Loj5xHN8XVk2oKJNBsK/PmCU+
paQb4/+Xd3xbvrFLgscMgCh4qeJTvJFfH/NsedM/NntVlPtYOGTa4UbD3xs5hHz0TfsReG9JVA3Q
cCuo/sdzc/HHt2qlGTNI1NznUFaqfb7BeOW2jHeEZFnx/d1Em9Eb855Z10coq8Me8Yi1h4xx5Vzg
6kZCyEpFkYfng+Se+Vm1Y4CzZoNDWeMDhd0Wo5jFRZuYRYjceFGdooRMaiYOv2/2VxA2ImsL52h1
aLr01Ag9JC2PTQSiF1PFFtZcY7txS6Nfp6jiInyyAg5al/yPwCo2gzs5RHWTSEnn3fJ6WAy5XGi2
DA1wBSQUReS2wgjIYzpp/+HRzlXyytV3w91jGakDtKalyfLLUQprfRtSFoSNdo+NHTL3j9HlCS6z
Ar8vf5KuGEmdy6dRU7tI2VtfM/dcAG9VlU/rkM4o+OGJHc1TRYaRrheMVZJojRc9holHv0cDZ/AH
wAMGgd7F2A9DaiMpgHVAHTMIc2DSJBWWuLY60meXTCVjB7TSo72PWQ3KDTypSfNz9s9bS2plJRh4
B+a4NDbgsxqDY71fNjuijt4Ugh68X5vrlXmw6lPKL6IawBYvYb2BXHGME1OfPM+8vT0Uz1sfPlkF
NopGHDEIOMj8sOX8l3KXrbz/vwmD9DEcLkxQ4GqAjC9u2GJlDyVyJ2bD3zAvA26LD3MnOlQ/dSC4
buDrt2m2KNzxUDan8kFpC306pmuj5ScxOZzpQ8OJfggvEMQHel8D607gwroQzs2LiOFJCAjGO+3p
ZVWSqMLhOk/Q8zA4uIepoh7E/bneP4Q6cJh1XErNLCahDbHZL908x0rnUhqQwW1cX6XpSrGpiRv0
XQ+Ryftw8cDVXU7F1jQbVNtIEgeAJZkf5JiB1NAXYsxe8Vd5sIrUmgJr9np6Q1xWLyYfDUbGZKXW
GjnqBWv/JCT6IHF3MKy/z/HyFuKNEIv156Bv+l75JoD0R2qbrTOGqgiEuJcJ7jYBsjXmkHXRiRtJ
3k2n50qWBZXpaVB2aaIpOltqwj4QiIvSVcG7ErY/4WBhuGmy0nYW77qh0ud6ACB761CnSa0WHeAJ
WOK/j+B276B8sezwCKiUNk+3dItYynK6EyROFjdlF5a/9gyAw1xSLKZ+44lUnRHUr/w9LWcHcnLw
MB8mP930DLmuiJHt9eP6hkJ1OEguDLxIJPQpZoRGj8f4W5IfQbFwekv01u6MM+tki+JKGU5y1OrV
qCSsWSU170RmmQ6kaRBhtwo5okNA/mrjTeLAbW3PjqeYAhEetFcWQJpvVkrGwziNdx0z0F5KOWrY
sHXlAzj34vbC6TmfLFHL10t0bneQpsNIBUUBVNGq3Hu7ctlVIY7tP99RUKb2wmjBGIBqTNFGOYL1
pZraikOKGpS3OmCXP/nX1JvgVRrJaV5KXeJN7OntX26RJDJUEQMO0hfEoxwoTDKczPm+bK08WTlh
Vj32Ou4Xn5/QkCV9M9+iLS4+LwcUzDSUDZZzsyCZ7J60VrSWhRAQtbTOa6AXUV81T7kd0rkWdWet
IKkyYEu7b+AzVNzC7HXv4hHkNOnQqLeRAb8oGudBDJwetPI+XKqho7TzOhywzz17v9mV/cGERz4n
TY4F+jQ2al5pvYCOYjgnrZqEyr1qVuhR0fsX0kKO4rJ11bRUO6QG1wNeqj6B9NCCQLvOLS+WD9ee
LPhOZ57PgZ/xWM5P1zc/mrG0Z2oXzJ4g6IGzSiNVCAMKZVFmqf62N3euuDYDuWQMxhylenZAI37C
TKMl117hyIIqo6ot7m8znQOkd+GgLM3PFpCkKM1seSS457k2BOE+HPC+sUXabS/47OeFlNaA9yQ3
XAHvQGhgmo9x/ZqH4krQz9gtgLR9IjnU3m2wVZ1VUEpGquFaBZ3QTSmmihAZvGtZkS1VqpDSO3lg
AZAdNInf0R478+SZzcD3H5MM9Nkz+l78DyZGQpOMOz7znpFsUzTH7HzO/8MqHeWjnNSwrOPMQ3Ru
j+R+WiTdczs7eoIsuKnUxlhT0d8vscf4Jzkb6V74XzvJ5zuMT0J7lc1gSuXQvI751vFDyyB6iIC2
irJHiSk2yMT1E2j1Y+Yidutp8YwpKTiHcuylogHjspQc4Qddwu/zemhWzdHTYulu+Z5GMnaCpbuP
Gz9GnN5+Ziyt9MGdoO6mibH++tm/wWJ6KKrCCEgam9MGKsCC4K1uk4vVCTtr8hO7bUvuViC3emEU
0os6dNE9EaAdCRTJbcuFgjiaXz8Nhp8pC1KPc80dTOws37fDbNbTZWrw6HUX1beF927kI2n6Jfn1
cWWKei6UO2zP3M73Uj+XKJAvtDyHC+nCtqNn6wdwq6dQ0RDcDGI77QbCqLBCdEHpX6N1N6MRitoL
plUXsg9eA599mga+NyWQvs1vVrs7jrjQam6kz6ZzBIQLop58orBRYWuyXRlM2/79aRv5Sb2Bw0XJ
77YCXSDc2bBONnsVpTCNcflzql63QIPmIlGLoqbgxdAUW2s4iMHIkiwOTNULvQ0ewwQEO85/vBZg
Gv6gcvThc8VQF69spZ3y9ppXThCHuiS9EnsbAQv8o+no2YpkQAUwUh7XExQ+FQZWMVmmFV5mAAQv
E9uk8B3c4G/g5R/bDBvxmeWXbvdFo05arU+eC+dBUj54EAPJshYKgSgf37LM6t0PjrtmEhLvt43k
QmBFF3wfVlBbpeZNqFWmlBMdiWjudZPiwCVUc1KxgLF5alyHRdpTm6aTrTZMLSzNRZi1RymwWQeF
Z1Arv9ARNn8SFY1SwCgmIyG2fcYVpwal01Nig0ZuNfZ59GyE9x13HbDdcZTFE2SjppAFiw0WOoss
LYlNAj147GpCqfoeUOmApZosSyzzRuu49BPsjNGGViRjVb6ApMVbMsDv8dygI8DuE+nX3umAY+LB
8T3NVLCfV+Gb5PYsO9E1DCcC6BoW0F//kFy9KIv6Oju5re88U5IDbL14SFc/yVzHar9f2x7kwhUw
GFYkLl6tU7yOfFS0dSCSs8yGGGTfelbpu9hySgHpTyqqIY3TukdFRGszkcBzcFX2ex3N/1RDvJo0
DpfPMAeGr1JiTorrGODr6aKR/xCCbu1w2ItrqcDfYE/q7RVnV0twvsfM0g+6et70KijGaK6EOKld
yIM0RaK53kThOjzTPSrJhuUhKCZUgatzAf3YcUpxr8PDIM83gIwfGJGa36iWlbHnlHt0bJ6fP7GU
B+KDWrxOrEx7HqZ1uwentLjBMUjAq81IJGPiw55bCIVglaruQqDxUXLxL7XnxmfBM8dyyfHQO84x
eDegGYphW3FMBqD8K6otEKtoFt+8nsQkEb+mMfH4IBzH/9ezbupF4homEzdMI8JoJ97bN/sDjz1h
ltagskPdaNiMJ6/xmxTUmWnRQJtuHp76Ilx//M7UJOXCh+uoDz9gCn2n8hP7oAhG5suws3Qjt0Ig
YsPY7E8dUib3rzKIv7p01C34owN1YSHFzs1yK2HlrOt5A+3KfDgl6oDxuqAkEwV59BFz+RzEFxoc
XANv0lR3s8D5IiJbuGJ3eBKomx5QwWubEcxGuqO1Iuu87UK4iB2MKD+7V59hg2QcCEpxTQoQARYH
AERShQOKcC9vo6LCTlIGemvpPIDdMpR8NXWuHVJAFKjxbyKuROSJHgoqvTNxIMIzLbbCWYYoY9lF
yzC9Bze6Z8rLNRJJDEy5evKOjni4AhNGJhk1qTj3i5hbVX77BmG8vGBsYPC9mdVzVdqjs6cilik7
Mc9TsWMkycX2K6dtnb6yR7QlkBnK884IXvfGt8r35VtZqm1jXmx/XqL957IjS+Q9Pbk+BuwPACuh
igxqo4i0B1zt6G7YoDF4T96gJBT7WwHseCyMoiIfUoAAIkQaQ0gFlIusHOtXZ/Z6k7HinSaBc1By
AuAyGPh0vZl73ajpPS25R2bsS0CbDn1sSGMivkbdbT/GHWMlofbn34mJCh+aSpa6zCSWE54+0Yga
jDDjYzQo6Nz+DqZQoc2lM+7S/wiYFqcQn0mtsdfz0iu++oZ+yZK9SUVw0teksA/wSDtt5wX5dG4V
v9Y72uaugq1u8T/+Vn9yzNNGEQAFaumlr0p4+Hldm7a1BUr2aPyH/0PWKcXNzwsfVvxXZQpO6c0n
DZU13OUSG7O22lpgeJKGAZdlBxdD7S1YKeMqBz1svnuPexkiNJPYuiDuF33yN8hykcqvNtrC7pp1
NhCKz+WSGCoNF6uEM1Fe+YIzcS0cyQFbZnMKExPOM9sLc4p+JeH5AJlA7cZnQxwTw/ZMT+yBHEYm
/1Z5LtVDLFj1urv8cd1vlmwI2ywNeb47LOgEPZ/9j4ar6FoAKiqxw353SLNW+kb6GuO6l5F2mrmI
HLrCsbD2mJI4K2ethkbOCehOhKeK17EJdt7q1jkhbgQxmYQrKqiSYmq3ZTEvGxiKihwP/hlYlFAy
kRZOLVrjOiTdvTEb4Cvc1FFhpsy4v8pHutZyhLBkAEFZFCK5eWnoE7DnBAPna+8Y97eJIKW86Kte
caVK9+U38ey/xUgmuNlWUXgewj5K/Rkz87jaI8kOgARnLn9fr0OcxTn7WivULihGioeO+lbwjBz1
e3VvwRnCxerN+S55QuZJE+y+hZeoQObZMHx6vKNNU5tZUbMQbxAG0JQL7uTcnIhTZRtpSw0D7qOA
3vJ5ONJ83KmfNCwngRFkZNJXr1Fmbu3DvAaC+Ni06gkZddde5rQIbTdTqkDTi+TXtReefKLuJ/00
HvmWy1GIBQZod3CcrqUVZ9xgraINT2C0pDu60EMI6J3PX716m51YnmKNbbdXrv1MdELmPvSwoUER
NChEGG8hgAR+PWISdqc3vZGMX5eUZeSbqN0RA8ObtqufyTCErdKIsQ8ZagbvW7YM7NsHdz5awn0P
deYr6t5Q+TfdJMHry43vLzKtTdV48az/xs7vzySB/IpUizPf4KuJffLZUBHO2eCYL6AecZabGout
6iBRXXRiUHTMLpfyh7uv4koZQ5JX4DWQn7vFDumYAQMHBIhVZ+7ZELI8LMiBXq3gVWEAhG5Ro3JZ
bNV6t8VdviTcs+rQq9O8n/t9rHPgXSWlk1y9IWl5nMZ3PunUhxTmfF1xN4uwWe+tP+v3wxBYMMyL
2pYhgBSRakrqnoTQ/DdI6eFfbYLGN/53/3wc03ZeG23nmo6iSq14G9GiJnLfWFie7EneE4rtvJRP
/t1X7yiC3gm7s72iOpXfaxhq5ZHXG17vgb2x3ws2qy80Uiwv4139gyZRgWkmy7YdK0QXqhWjBqeK
DXyHTBPTY9VlNGZFk1fO6Q9A5bcVzHedLkH1+umqwiTDr5DIGNncbriwAVM3QEspMOjiOXkawOid
sC7WEdk/wMBvTMcXHb/hPSu3eGgabfNugJ3DjEneFS6XMgYzy6GImEYU8lOf3S2MqU3F7+PaEvMh
qnSti3Als/OxYT4XFHHkH7ClwwkzJkXOTdQ305ElJ3eB5Vqt6J6E7PIfZiuZsXGuGk/cxsv11P0j
3oshKODj+M1Wpt+krhGvLnddgjuHhWZRuZXhM7Fpp196jITiOVXTXJpfDeqeKHF2nUM9puOJS3p0
r2so1MX5FoCljvkG/uiQjKQflrOdz8beBZ1b4+FuYfZeMtgPZtESRFbdoLw9JJ6xZNhuxdY7D3LU
qTSPbq2ZFuv/c+Ybc/8iXZ84F8mVtoVEXr97RqIbkDMbozQfq/zqg9+IxXl2x4/DHM0hRDKZEsKM
S+oyWD1nkmtss1ibF8QOksAWeuA1Pzt26DHcn3yHALPB/QsxD3/sP1xbExKYAOs1BvTNIBpfCwu9
SOLhJLG+rMwzgyVYTTpLT69NiAVG72Hjzeli88d64tFE44fArDDj/PE8oGG3XSKESAE55FQd6GVX
f8jml3hPeFCq3C1lTjzxBXlQSySzonIDUjrLV4ANLH8kgUR6OgsJWgOtSG/R/AjdAGNXSFUHwqDF
XhQO9M0QaT20ON4NFLZQAQFTC+qpMRjWhe1RtSfMQVTuZwkOzgyaDrvOGY7TMdWnSgGSgWI6K6W4
y3vMBp3quQ1fG3qcpm7S43V7W/AwQDWbCcnHnH3040zepEetB0dWYwsfv/mCUnuARlPisnrG8aQL
pyB69JY/u0Si5KxU2TEevdP8Gp0H3eYXx1vs7y0IuwH1Ypub2wZIyk3+svxci345z623z6+jS39N
heTBwbQusDLXPSczQLHiVIJBRYmgbW0xOZHoBg3XBh41HBJOmmDmDnckfoKojVUyLi9YsMJWMTm1
4Y1zWi+jAj7IN8x5OS3nnBI7taDnityaJhLjmQ/w7MwuNsWxJUhcfaqrIop+eyS5Sw0zzoMciUql
RfWgIS71WI6wWKtT/TCYnImNPIpsN2F79ke69WA2aDQPMvRw56fvchC1cldyUR8o4S5pdjxtT/v9
6qX0Ems7huMADwgONW1NuEC0AJOOcEjOzYzbLOHD5C9oIHl7O/YDuNA6d7ofZM8acMljV0ZxLFO8
fsKye1RUAgCKifaIjHuaLeab7QG8y0GykJetuaQOxYQ4SgcPb0f4yEVpUpSr1LWAT6QW9T7kwwjo
d4hqo9ZL4Vufu39PsXE7m4jomRishqVB7KSosm0FxxQJAo6zOzSSm2/4U1FTotc5c0iQYVGcgBG+
DJxOBrhW9NFMgPHdzwcCYZz0czOZGeoFCL+cievrRVL0KER5EJdgiFDlQOJt/i5MhOIMO2PVy2Mv
ZNQHyYSVNDdcld58YT0OXRLFcC3cnER5fHSJ+pIq5JjxQzIZybtg6qWlLuPDzCaPUz7p5xHIlYmE
4KFwTK+MsMNmtyNKSSFtAvxRBOywiYVUGUSZH+lYeUEK9KAZUd6mbaFkEgYIKeMtb9yfROC+dOFH
yFUvk1mK/PpccO9vpuYdmQlAuX/O7XhdINDwgN+HPkmueYnQeZMkyimFyiLdoTEaHZUQvfuKbir4
KzIWtJRlOuu/YP5/JJjUUWZqNREAZYZVoklNuV2gfkFyEGgU0xn7iVD2z7j01+z5ubGiBAOzCgzv
56YOwxBINjrke9BKu73f+zPkVllsWCRs13q0QwMkx+D4n8Hsr6gsSkqZxBOeulpLGXNsiRe1tnx/
LYarvnK0IEmyclBTA7L6ejV8hb0DgzDx8DYOgm/HF/p7rxAcPyTeuRN46nrcnHNYFZkWIRvgvrd4
Ed7YKXu79MFWrzQVuj1qUescuPYJSYMFL78iwywO/dK2rTNCe2oxaHMyvA80X6IqTEfnyuVVp8st
EYJdasF8VJ1m4vfn5hqBRLi9ILbpygjJsL9Gqp2+YlY/MYlHv6m4Wsa7+LMYctI72uIH9dnPl/uU
VRxqjDjm3Cr/Fglvb73eotRxtzQIX6Eak0zkICdOcJdGDxVCXxH/KWWV42z1C3Sr0PkgSNzTQx3v
1pFSQHHZwtkqMqONfuBJmABaJ7CytnVa/pHcRL3FPqfNCHByh1O3bh3aWK7lKdjGVOupEvO1t9Xi
pFnzDPbZSrSRYApTk/OmDdytmCuDMAqTaZD+HlpaVM6iqCSlliRKXNb9mPI7/0jYLDUZaW1KPF6O
IxlB5MdwKq7PzCfQyzUXaDptJx8tFJB1ASxcw7i9cVDmpXmJSwvQZ7i9szYieXysZ3ALaZPmkysP
q899DBUUwPWnU95N9adpi6YtjZg9hc3enWyThODW5zNZcTug9GHFYexeCWyWwhxF5Rcrykg8EYYE
Z0zKHPt4r16SNZF3LUIMhqlQ8X2jCe9JiiECDFNIq+lr1qFQcU2a6ky8ODo5MhPyvBM15u3aO5zy
qgSHPUrsk2hlFCBcX7eUHhdszZWMLJXwwSrYpG4lqwPCk5CQj7Y2otgAM+yrR367YBUzxTSWtMGM
Wt7AghlD2cklPkZ2JMKz0FNFWd17eplev5R7K9KxLLTDqI7CpWIiP5J3+uBawzf4kIVhHtWJMgGt
9a32p6Cmta/kRV8j+7BzxGXS5BJjZq2InwIHRnuvOSszsZWgY7Ul7JCHanY2YJh8Rp9JE0/6cP6i
WE/KfTwW0Ilerc1rP36Z7uty1s4J3gqGIM1v22NmS9MHuE15tj2Z9NIXhYFZICB8ITAIvmkbp1+5
paKpy0E+Av0Z1nQlI7lS6kgzNrSdAK3ZpCd2pLMnc6u6W3KF/B+sWWkFoQ96I5aTOoXuJ/80D1/B
r/g1i+v0GA9izcKmXR9i1bynYN3nKhBLIqXOH79HGA1Yo6H8xbTPUJ+/HJKyQQaOII1gjiUc6M+5
eVjo1UlZfRecl2AVEXrGbmpxU6ExOewOG1Jfdj3F7dTQ1+V2qtp/mm6x1hpAeta6+KPyyThB/lqZ
jZQ+lkKXQ1/7rRi7WTs+UWEZp2a9BBqechO3dmJnIEPkKSGc77kIwt1MqiX9CZw3qSPz2qp90caG
v6RtNxWUzvZXSLbUsYXMUTw746XTkMqH5AGdcYYM/efvh62ZzXf9fRIpVGt6+njqrRmtcjPv65PA
U2Ds69tmT0nguffHePZc/di9Z56U0b0ABocGzuoKIUrGhAS7YWpNG7xOn6tqBysr0/YXImdmHF4R
99g4lpoLkOz2xATskf4zC522NezuNy+7SHZzOqlwclylNx4QDpSgzia7WPcHKewmaEBGcqqh7JCX
Mkq2TycSIU9O+3XK8/B7JJwWpcIpKSK4leyO98v06pDAhV95LXaR6m1lazGlwWkGUvlxGO+Hlqzm
wcb46e46e9eJGP6cE0SFim0OnB4nlrly2nkyAP58uURw9U20QqCVYZCCUT9eevv0pPYt37fZ4mIR
+W37gKsbZ0Vy/MgYqKoGt2q8AfzIEQ1jo8I4C0N4WHy+ycg9x+Snh60ISM8dg54Kq8cxMcZkfokB
eyuM9YbfwdhsS1ruStlqEbvR62/QL3E2cmomx9wGXA+CpxxN0tuw/y7DhpN1vFkMQN8uFNnn1UsH
sytOHNIPiAvkE7KegpCDniizvQ23CUREMgqmvQXSPhVN6kz4kTRd9KANtHh2ARHo5hqfkEDyaioK
jkyvxDwPIQjfz+0FoSsEXdANTt+Qsz2VTij/crD1UFikLtpuoG9tRY8HRZoZV2tpiy4O1NBbSexT
cWqWYGMlXvJholPsS/VCMdtvlcyDQ55l5fy0emCVIfYvf9lK2tAZlNP5enPhOIQqBOu3B+faVf3w
sjHwEKTptcSVLkkhwP7GWkOrEUoqIGhJ8IqAEBPFG5EF393QXVrT0GU63ggL1XjhUqVWSdalvBqo
AezNplo1e5E6p3N+M572pTyYc6N672f47yyKmelPhb6oQAWMWorfRAUwQqOHM28gEvW7pM+yHPDD
+4319tl3zFDrKQW2d/vdrc/FQNXgpja66a0TvMDMsqPUf69FEIklrZAVDwomHJH8IYV2cARJfdjE
iyU9KSI62pipmkma90zHsAnlPUvyIJag2sg5Wn1p8jDliRMnj01DN74EG1x4L+YfNMviZLUsxEP+
r6fKXk06bb4HjmENEDzTBSIw3867UiH98nWnbMcqDlhji0qPewRPXUlyJQhPNnLKWaF87R8tX5B2
RkWXelZVxcj8fvDrzgoNPaBp5RsibF40hZcAb3z4UWkvLGhmXc0z2om4T1tXlPChZlFwgubK+2bJ
44G/UlOhzQvVJ3Y+Kdm7jkUYstrwQ+bowFgsJAkGKGgpZuR6dx4OPV4jVvboc2/zXrfVnCS4ogJd
/hRkUtINJwLfz9PQtlAj+XrcY/LhZdhnLaSpWk9OQkYcrVxnf3aRgbaUfuE9ZNMEt0gvCB3cltE4
Ykzze+qAAXL5K8ORYLcliMnMP+0cxHGPoBuiDiTnGZRh5uBsBlOdNFJi09DZZb7de1Ey8+7dVDek
QNO2WbKvYk49OYDRbkSF5ZgXy6Zb/Ab8UDInsp8bdhDWT1U/o0N3XROxRYHb110HVq0fxKmRlYMz
yANW+Zo5Eerob7VZiuFqb9aEiiQEBvo5hTrJ7Xjm3PUz5cx4oRA+rP5YB6E3abWHbB6w1JCCoq0R
jNfpIhgdN2J6PV6KfLqoT2Fv5EZ3ubY5+PZ+OniZRQb5drt3hJNvfHctS7xBdhbEZEHZ25KL12KG
7npQEEtU8SitnCLhkI+jKKOgHYVbHU1bG3Rxhap2y0CoaPygT4J6q8EAtH/7V6sarBknMqAI6cHJ
Dlt4X+NUR11vTV9gjg4EkzLxlpnPGy0/nH9v/bauw/KrpQmMXauMZdleJxGJuS2B6DnFANwatINY
kxpx08gCB9FsNStEmKpsVRHjfnd2z2M2ky/MMM48nBbB0GN9e4g5o5h9V9CNvIHgLj+7fylZyF2Q
NyaH8YJIiMxXO1eP8hykrDuQRdCd8P4EMS8yKUMnlpV6Od58NTUcs51ldK7S/wLz6KNZ3PcTHCSZ
KI+E4/0to17idzC6LuacHnmL2eGlWFbgvDOMvhrblfGUTUD0cDwCnIV1hqgVIOqXDLt1KvnMD2WB
icmEuLY6UzRkgoRyWXuVFpEDCqRV3al9dj6/qM7T/kfLkRj4i3Tn54XrDmIYL46PJztfLXP19cfC
GNgBTwim9mSfXqMI0m/RqkcDDy3IWvW2PbjfPYFD0rw6Orp5yV/bg6aMevaKN9uFBtU0e+t4Wj7V
eW7rEKusvVFW4Ow6xK7GST1xtzFgjlDh7G4xaQy2Y4MoC7KV1r3XNSmLahVL9g66ir1moY0Usz9V
4xu9LDzfN6zDRr14dRBSXMsttyg+NlsikM89VSY4sX7ZbehCSxgiYjXFdIXDGfUjbzWu6dWb9LIn
VIzXoYMAP6w4WT+HNBzAI1+Gx58BUjMA0GkdJGSVOQttsOEPBdADPtdBA107yffZOUsX3gkj7GJt
5fFOJLyM9Tdu23/5nFXMrNI29Xl1pVNuriycQvvaA+k91V9GFQehI7p7pqbrurZg8hsReUI7ipW1
P86TyjzOMuKQjlTUZrakjEkWI+7vaevTxNI2N8EGonLJEOjRLy8aUZhBBwmL9Oz57se27thCUeNc
nuMyQFKmWfL89BDyvEcHaV8npngusOjpy0DNlsMotV9fKXOqpThNavud0n/nJUFEUK072oCHQAFn
7gnHgFIXp/ig+M8m90BaY2faxaposydjAa1geYxTMmuOnl/LN4Wz9RqLGmjmtxnvHSWF0HCqOc3Y
X4u0VABVDtTj11z8Yo10XXUgDWii0vXlF7lGSOkQInPSVUmtSAhGZcT6qmaeVDCEEFojTJhvU+cq
XefGvOkYyLAlQSyoNfeiX9nyCU48tN1mQHVFlNj9/0p7W7IgHQcY2oj48f9ZKbiRGYl7YEefGcsc
FtqeTN3OpGl+SZeLLnvCMnUn0Gk/V2qaKhlUCvySt4G6lmrwzN0VX3SInNGTLcxMyCmzSErmIMX1
jrwXDfxSBmHgnzLTdnVRqwQ+2U5AgAzuM5MWWwLnXlIjjEjV9ZSob7p8noRDAhIAvitqkb7qHiut
lyxNFzamYAfDQEzyg12kM8h9G937j64COrRm7/nghu4rYCWJEY/ZiL+ukSyJ0uvuk7ZkkDWeDj9B
7Bu22DjZTOD3icgFbdfkWxknE1GHTTyM1zG5NEOpOBNgsTPLpNdc40U+7p1550W3xRI6U5ffAEnY
wi84xEIeFMJUeO7iFpGTzHkSDExvsFncXv8DeFJ6VRTezkalAHtLmVZAXXSzGF3xCyBYS1QnlRPT
xmPzh2YruSMDPBSf2HwnV95Tm9zZQr5NjtJt4m56YkwlDfXR1yFscga9K8hfKp9O00QzwjWXdenh
SbkhnUdv9XIkwgIX83SRIsUk5pZ6tDq6hCCAYVFwTNVBxxDqH3C4xBTf8elIA9FPEIs3/TC9ma3u
NSs3vJAWYhfBsWS3yRukE9yVA5Uhkqfc9PKfwgmjzc1USgmx/QCJ+84It3VR4w7YYPdZR3TV/PbS
9e3bJ0YWp5wd1stZYkLZKj7N5T18Dq223lhZsqd/4X++3blkYNCJ++UYt0cUDGGAFS2F+OvwTXco
zk7smt24lslVjWA8K97nOyEs/qRhBnybuxQN8wiDzAB2ZSk+oGuMo6JlhmL/q5I7L8FWJSNWzElm
LQJwSCtTnjFVKCmxSVxdb29Y8OkSY6pxHif5zJ6yeSeI43XFSDQqGEDzV8hYmPwU6zaKhtDV6us2
OlQGDH2nBjpgubkpH5RRx6h18cGuP6JSFWF2vLU35029/8CclT+HvCKCwM4t3hWOn12rW1H9fZ28
3vuss2m159nmccDMNOOYwkdC8TkWrbJA8tC0eeMea4LyyikfVmpZinViWfJAzRb/ZC5y+7aGHNnX
fUzQ0QrJNZAr6a0phyB0PkMC2VQF+eQHv7oyJG2+rWlG07kSy1okKioe2FTtbSIAa/z+WNRblsaJ
9c4J/oPt+gFQ7QKvdAn8c3MX9IYMynDtP+aAl2WMwz7GslHIYv85g9wHRtnSXMDehZnTUlpXDEbQ
v5cUNsHTqPQprPrmCJc6gNpoBtWiN7HzM0Oca17j3e3lkYvFK/4dwZuuh5HePvxumAW0eYX7Bxg3
Nc5QZaOcTP2HZ6Th6VWXw4E6s+kMQv1mEdZkaKMZGYqKJnGAaQB6lFUcIH+C1fhSrFdArx2UN5Kp
qVyAEPkLzF3jbIGjnfIoZMPDwVDJfnAoduX0BpN6gDsk88qXM6OZtWGmd2Mo7OehtAar6aU5Pfmb
HVI6OabFWFkFCYAEiwB/uhRBuP+yyxu271RBxsR7XJIaWSrn2zin4B/s6AFmchRULGKzrwL6l6ok
Ur+GQIzy+tL8/dIz2vpP+OCWFTBCpDVozfc6U011RSngt/5t88pPSfq+XWRDrl/6MVgCb9sYracT
ZtAp/6QWdMbPAruMaKjDg7/r4QZho5wCSCVKEUCllgD7vIxJgAIbbbTCuRN+2Eps5txnAiMcaB+J
ZQuj5Jxn1jhqxHLs7sh/u+zwWbz83wC19CB53JO2BxMrAaj+zcqHYOf1F5rahLow3nn7Zh9BkBTW
Dnal5mtikluFPYOzmERXxWq4rBvo5V79ZyAFnHrFJzgdxAsBaHVvDFfrEPGJre4qcDbiukreYizB
AtvovkJellQvKpQkkrin1Ti1OKXssUe65edoNI1qXOKR2+rVC0OquJDCsR4Mi2TultMdPBsipK/b
lCP47hSh6nprftCsY36uFr5zFotllwfOn43PyUG3heohDzKyOWUU2mqTuBvGGvTM22ObX0QIDmOH
LjeMGmFP3GRT+WAJXV7NX1guvdeVA+YO/hetSsIMnlTgp8NbzGjzKN5NIejUK5AJVA9rW5RHncol
EkUzkUDInFQ1hZ0wR6ozA8eJ41QdmtuILSM7dbj9GeMZSTScl+n+3BImUwe9nTQGhU98VXL7+cS1
1mgjC2VJlWPBwoE91LZE9QqQyC1JmqR1dWaRC0ck1bZIBWz64VtEVD2GLnhtiheMUxNHSNv2gMfT
D6fJZbPEK02jJp73D4jHiLCBzOLs9kk9imQnILMIUBwTkFibwksURtV3xaO8Ik+NLNaa8aYUqGrY
cOZmvygK5UbyebwAB46howoZN2+gg4qkl37pPgphccsK8fwP/CLqP8QAPA1z+f6FypgwREjDCKqY
5LtazEP5biK+i9sW09YjyzQFSHwznAnHRCO4XLJSGOG/IVor4M7oFVVX6WRCtTnotvoJ9pvA9hQs
vxO0oE5P6WwMF7lkeaHW7pY/17t5Z0sHdOeo1vuOQEC/kYhbTdeBZNRvMsY13f4+EfUKr66L/53E
JGmiJV2YjoRsjMUfZe970dk6WrBJ5r0FKFPLknnHLFH1nisn8N1TlbRO0Qy2wAHhInYhcWOKQ73p
7K6y+ual3kd/csdFDGx9Ucd5MY3oBZaRGG1X/Or8G8oQz5V+qWpVBFTI/ZH0nJvXjko9AGb2pyfr
A6FDX2KSdDtSnI7d5U1+m+QYSrrhlYqMo68zMHdl7biZyaBw6esM+Ff3S5FkxpevC8+Z8fkILlug
TB/qIPIwkI0ze39cVgWKtZhU3qem+jEm8txYxml0GXQe6GEEAxwF8Yr6XDeq9BlaQuKcsxBiu/NA
rCZk42reQMQjflBod0SEqr4Puka5BZPw6zH99CcZPgKP5r1BOiGbJzfwWgId28znKpsB4/I5+pL+
2lMUz7eqi3nU9BHdEd8JsbziNaVIzog3exwZlqaB+wQ9VM0/Uu0B+8zBwVa3VtVfiS4HuTSTwXt+
o8NLr41qIMON5EM2u1l+jNzx6fYdecoR5T68h02ya54p7yGPsFQknvJgSK/WKf8Z1ZRtB1yQCyFZ
VEGIwvqWxSEXbC2m7EC3RDflDQm1aRuQmaGw1pM45ITknu6n/bnmXVAbOEHH0BR8zOW/q+LbNZ5Y
RS/WkFNyPhsZtM8uz9oLUdxFFVRCbDDmzrIFW9LeIJdQbKa6zUhkRwEP3K4qiDm5L+GQK81pfJW/
T95Klyg+vnVnGOumjpAPS3NmJyqS/kF9Xi8faceyYXmtcqmhJsaOpV8pJdcDmL0WUM1q9LGk+7Hr
9gitjgZgv8NNynMlhmcHuR9oGz7xSSY28kKxG4fGjA0x2XDR4K5RRrjB6p2gBa8CHuIFbv5fYVk9
7utedl59kBxl8Rr7Te2OoXYbjXRf2MOYf77yJ6yDcRSTZCbZysivK6jOM16PO/Zr2W7qPmqoV5pW
t3z7BgcZo9wGQ3p2wR4CIyCNnrMcwS4iUxMqYTVt7Xs1Fp5MUX1O6U3YSB5zG5O8xoaN3r8nbbu4
ZKBvSQM7hiPlIuJNPshJsw8uoLelNw2Rkv9qLyKZbuzmS8Om/6c/F5hjcbnFXm/5iwRIXYmojgII
ZVpptBwV9Iug2FZreAD6bN7jTsv0PJ8I46kUV4rlScj59XIpIC3xdTTv4rFyNMgaZHTJ0M5eoYVa
1jM8LKZkNAApYNd0hr8zUzZ7gHEgB2p5aITuR1L8m/VbuIIzCHlSogcNOYj1Fy8n06IE+bnKU4dX
o6w2xN/nhGLOQuQ8YsHmRjSV3kWXtjqE9uoVWBigHOKs6Quds07uLTFwXHYnCHHz7hIW3O3+jro3
5zLrABG6x2RCIcYxGrBJPFzheLABNg/LSor9d5GfNDMDZXxEehU+ixcrUahhKsR4yWgdzxbzrsW6
ES2AV05sANP7es63ygx6Ul9NpB1Hp3nTfYeskvUbhVuOXbcAdt9wn1eAIR4GujKe8rdGUgw7aAIn
gwyYy6UJ608vyGM+zrB9N7I/rIXmw3JpPcMUnpTHrwixc9yuUHH/T/hyt+F36nnEDG4Vbj6C5d6f
s/zN3HkwoJ8CQYIubQEcEtFJTR1LiN3dOjTcpoLXisHiaq4xiQdMVL4bgTBuxzkw4JKGFRGjk4ZW
aebctqfj/eS4B2266ex8XGmqjFJ7EtGx3AT6PVJCe91NBvSU/h2bN762NyxD7zLgmQylGbWULEvt
hVBPRzBjjyXrCxle5kVJQIOlDOvI/hBSHxigW88+sos4XfQqJkxz7fMo6iCq+vow3DxT6JefhGNG
RON72ZuTLYaW7jR8+9dEWFQzLGewo2tljmgOV6qY/PiQPxybBiNY7NOS9gMBe2MZrlLIT1nIKrN7
Uw9+OgCSP3IkQ9fPo73cuu3QxWm73D4LjU/hvWd1J/RF/hQQYht5aI7WqitkzpSFjLx4I51naTeL
s3AU5H32ZX1Bf3HjSyOQwA3YQEse5UTJE20ZtoSD6z9Oen4Tmiy03TM+Kow8nGQgEVjES/vrA0IP
Cbkr4BJCjOJGiHKGd4Yq3VZ5/vJurtcoNGX7G3KTEYMgNelbXkWOSLtGgVtRIBoEq2fWi0TmbSG3
lJMsbD5i/VJRKjouYvoHHdGfNpPzLvewKbqPi11CAzxN80Sucs0eKUR/vWFrqUwyWSvsTpo3IU1F
5ndMpqY3DS6wMg+tgV0Sr1MpJgHeWK2IoV0es3I6jpEWVS9UT8AjM25tDniOqsN3+D0b+L5outpF
1E8Gs2I7SiKCwaUI1kQbdD1JDt0g1Er6k3QoCj6MyyV1UX2D33d4WFTma82AaNJt3NTEtauTgoDO
rtkl0tGtZ4NAOj63Xlcujg/4ZRyttf1p84CAv1AIv80JtPjdsdv9L7e9eGblz+oLQhd2mLL5L0cL
AqD45UYysRKgM2YxqZCmZ/hXawcq5aZ+n/IAtWFWQt7TG/xxSrQBr6A8GgDflnhsjiu19oYebcFr
cpw+pshp6qw3qDJCZWPogeBUwdgPIOWDEGJUK8+f0O7BBe6V8kis9ERsXV2BhNCp0ieHgTbwnUGO
YDbSMKWQ+y4S0HNDsb249gygT3/M/jjJF1SXLGfzgFP+zx5eZkadwATit32gGH4yqaMtRFBycqOs
RHQcFxtkDfA1ylvZNY4JJZgix1PjnYJ+qN5XF8WupzVtwpFAfRy1fJ6EalgMfjDdbml2K47Vwamv
v6dYXrx3pH9xRrWXr8D1G1375yfXOY4vrdW5/LBl+ROYtNolPvtE0OnAEfkU7L1lAfsW+M+ZTfDF
Er90TnsT7CnjmT35FlcJmK/Hq/AdPd6DTvTdbPWSwz9yHd5OauTvkuWv2fyZKosYJFhD5w3iQFeC
S7Mf0gzcclxZXo3sf+A3/6+jbiRSn4813RHg4+PcJPT2hkYx1LBRLk5qhgQlICyctisaqVSUm/AH
RzKFhaljZWxRx6aPFL8Yxy0UthPuvPBExbV71glKBKPGdHMZLRZM/agXi+y5FMYiYetK9EFJJiwz
dL3o9KxiMDfNSfCLlkeCSDcSM6XiS+QMFvYNRqKwID9jAPkMKFePhSrFvGi44Q9EGTJeCEqPKbp8
9jn7MSYXORqT3ma2M+Ax694IA3aw9jeTUHHy3gXTrFJxaTZV4jpNucJ2MKWIyu1gy0fiqmv/ALIj
/JFbNHzhjecgbEqxSunpRlEltd5npAYZNc66FcgI2hrs85aBslA1kUIMljxmeihoWugkRi7zuGS5
TKZjp6vJGptBkTGtKgNAzShEs+Db4B/V+kN4ZPNHcZohIxDx3oLE1ApUKuwecBFQnhNBU+2eEiYA
oOTOYPCYxt99BJ/RO10hACxGFjANn/JlYYHHFgmxeZZaLun7LC8dFadGXziUetMPKvbVONnqDbP/
XexROhm/MWL9xfy6Z8Vv2IEHWAL+eQU0rRi+U3lt0DqZUj6s9UI7UoM1W/hVfoQmF5k5pvbIyvQl
zLwvrrRXazwRenA0l620rNzvR05rvpqb0rxyZVAoSOnTWmH07NP3ExtSa8yPGJiDrhB+R1z1uQSH
yWaT24B/X9U06FwX05Kx8Tc5deHizP+khAryEeS0FxS3xEKIcxVl2obrMTITvMAhgGI8RQXvzyDE
KDzfCDvVB3EEf/G6LOGxhdXcF6I4aWk8SNCcmzlpvK1B+Iz7ZnRsxro7mDj9kZNRpnR7eMRwLB1n
V5fcXRwn++1Yrp746LDH73ddCz8Dv6scDUu5HvP3mQFQtjN/zvseJyfWg9sbafhSX+rvZfRNj35C
NeVOrRNwBTnVyVTM4gFLAVY+vWWBOhvUHpT44c0wP7bUdV4bmQONwCDTy6RtB48t2wtPFxeUYPnI
U8CnaVPacXPx8u3xRXwE+5n0nzBBXxvs96Ax750RobFbD4fLZTQHDnbLK3hBVDMn/mLItbk2oQtg
TWelrvYH7+5NGAzjs+++TULeKToGKdpfNQkT7CJUWkDBd4N3nRVOH0aSmyJqQpARzKkZRqwgq8XF
8tA08N9KsAa/bg3XnDfzy76P87xhmUX28OlRIWj2zA4COfiPIdvUOLnMvhmRXrs7KZSZS492F+g9
MV45Z+LiiiOc5pTRI9xi1Ui4IdzlhO4rEOSsPziVqH0sRk2gCYQZ5YVqRhiBDhz5sCaq3UPuvusI
DUuRGBh5uneU8odgVZ5R1sl3kc4Zx58duEmoJG7rg7etVJVhgi2J1BrJsQHOlor2MrbeAlgdtFRi
LInPKiQEOqtLQKuaPp2yMG5MUEkB+WRbeDoeJOjVstB/hT47G7OGMbfbxA+fO735e8M+Q2kOxBgv
43DWPJNASWO2jraRIN2EfcAhDMratauyni7afjaRNPKtJoq04vYxSPbsVPjW4tGQCjVABZ2RLoFp
MNzPF8oEpAtt4C7E7Ln7dXERlwt0VyR1r8hLNe8H9F538umdmMMY2RzCaae90/CGPuoZVBfO1jOO
BbnVO5TFnk3KMz5JPMbIJoTwgrDm6vU+pmb7ru8blWoTuAvqSwUoW2QQGptLqhTqnxkzLUjLWUS2
U6Hd/t19nRTZLe7WadKjg6xPVMvDWkQr+/OhBzhqB4FGZ5jRBHNDayB53B6OeHcsKseoriDvfg76
hrwfA/fF0Tzc3BrSNsQ5s63nj2TTkivZmHaF/sjWJg52vUvG9E6Z7yRKs1bcWaKQHI+NF/BJg9ip
10vrngZDpT+v30/2xHvqCUmv7zzuQUIuL6nHdPp7JXHwtEv18KDWxIWpBPQbxuEKfIjz1VLcHO3n
yooCShJ1VeGdSWJTtnAr3n59Sf3Th5iz8o7XF3+q+nlwgvNWeEgLFtdSP7qhzmaAXBoG5Lbqy76F
mDh+yB98xcvwjYau2iQHMRQ091VuP1+unWmwdLCaq7MO6+QQy95dXgrUO+PXhdnMHjb0Gw3UxHNf
7+tvFCOPLMKf8phPU8s8qcrnZExFYu2ef6pIXFokyFPdCopwIpSXYSOQSF0L9s1E8yfSihyxFYhw
X5MM5cbuGicxHlA8RZkq2kfUweVwvb3MrE/095Kn3xLGMwZlkkJkGWCi1TYCCaLm3u+3cUoTbofy
zt8g12Gdo4xFgWwS547mpHckScbqdsyNC5VFWclbANjR0MPjulOpll8/7pyTb13hI3KMpYBNVCxb
xoExgjjaydIC9J/LLN5OKB4wNlggoX33VL8iginh4Z/FfNIEieGLIDJg+PBsFZBt3zdy6kYt66KK
SdlhvwPRCwNyxdZ1NrkOxzRGEflUkWJRD8iVzXgklycy795yRCg7COcSDt6WwyU9Hee2q+ZCwNdy
Ml1R3cHRLU8kl5hnTYxY1w1fD2FaHd9taM1Ah3iPwVKsRwcIJaCZd8jXvtJJPkgHCSwYA1ZjE47p
IGM9caAba0GHqxsB2pRDgJU3Ii59XgqT7rZs/S5AfGcKZtrU8E0hcf0Tk5FbGkDcJkJD6qmsbwW7
DIFSPKThimG/iiCuyDrgVeA/K+u5Nv1GxcobwOMTU8mNH9TEtDuS5K/EtgfQh8CRsNwyj/zsEycl
Is1p88RHVtTy5M250mwK0+aHSKq9eTuMyY7EujS6XrXoFv2N3LCT6eIMRbT/8Oh48lCXtUDUEh/4
XJY8mpfJ/AoyssynUqSNKMiQlLYiyWg1bwFeHj15ijqu+G6zcJYk186rGzr6KvRbpAqERatg4RIz
f3rhc+v6mkNk/hibZoU5SUZBO+XU8d4aROIjUZlzrjbi9hgiUFSryoHnclf3SV55uorM05B4YdCW
C4cl6JbbbGTB8al1Q2Jdp2Le77N5My/r9I3D6v8sSAAf9XlrCoZw7/gkrUxm/xGW7RWdSXlsJ5l1
Re8++11uzOx2sKZm+18JAJeyVJZeVMwNGDIrZraGWxpcTWxt7AJrgw9KFEk7mY+8c9cdmMGPlhKx
1z1lcS1pjors8SSjNfglpotIlcXorI72OwPbDFINbYM1+XbBvS6F7NfMQSOIutiBuAFYQP6afri1
HUcx2HZtgwkMZUrGj/cOtZgM0DHboGChhltZ6qU7LIVmyYXb1P8fMRaTSyI29Wcx6imOJrVpRjM4
uIR1RvnyQiqxCVtUHKbmzBpgOyb0h0zPo3ENAbgfEyFPAn2iEUlKh1Lpx0A8CC3sPYP40hUqUl93
yHqsb7Nd5h2xzoqByu9uQKZcCOAwUTy9LS5/k2Y7M0chZbxSM9BNKUyfWwYc3JKFETxCkBtdYvdH
BQPHAHTzCPwblaleED5lqKsryZukXyuPQj9EsGI4SE+5kOmQn4EkuKASviEUVMMyLBto9af9QzgG
H35uHnCgWbQahQMwKdOHG17Jq8oDXsrHONQ73M7KDqAQlbfYyVDyMfaWbes6x5kxDZSOUtRmgVv4
u/XOV62DYP1CuUl/ofc6vRj0bcXYq2hep92z81oYFbRVs1T5/Z5iMeYVVGc58KLV7HPpA2PA5sEu
dQvytOyzKu7NwrDWxq7iSv7+Vm2JQdfT7n6FtIlwDXQ5dalmdQfR8rDRDCI5n1FH9H7O50Oq36au
Ma1RRsS+SmLYaRtHhgztGgXYWD9HTUgf0Hg4PgPdNN3O8Get/7M1B8Sy6f+m+VpEa2CqNcKWW64p
fU7DcedXlgA8Jcwv8yd0T3cb/mSK7QSzVfgShakpLyOKboYPkNxlO8AQ2OqV7Hxc0ynLv2V/KleG
BAYHL89MoU+bPBMokOhYzq7KkqyQ0GiZPiTyEGAr0oRYCnGtBArv4xwQMaUoOEIOtTQm4X+okd/c
hDEv2Esbk5DiT0wXs+uohzvbxIBJ75yyN5M1YsXz9cRGYuYpkLNZUTTpRk/rMuwwRBhUTyWyd5wT
XpAVT9JrotO93ZijMojUUMaL5cq5NM9/KqjkM0FjKvNU26s8ObK1oYXES5ZMbjb/5OC7nHyG8W9i
xNzBFemPx1AgIQR8MVartKDiUGVdE9sJDDBql55VEsDwHbBOc5M4055TZe/ET8v8iXyrLIfaaO1O
A+YaK52y4b9Wo65yXqD6scSdbYKMl73uWuL9GmuIKAittYh4MO3Ns2LkKu2kfi3uTi+9PG+adfgu
NGr0CjGD1uV1hb6JoHHS63yqFLxgLinxgM3O6hry3nwi0QXlWG9yPfLD9Xq2nakfzKLW82170FgX
gMmypNK+FUjDlW9SBda1h46fLrqyzUJ7LSFbZ3r5sEHxdQE+0BJqcItbnZ70b2SmhZIfu4rkekK8
L4rQ4Ux6xITM0xQpRsJR5H6U1xhGWsZA2wn0266oi8GTWhcwr/LyQPUbcyrEYpaZhprB+3lJ76Up
1AtS4qS67MvpAwTRMIYw/keoq/3g2uLjBQKFQNtEHxC8jgbeNct7XknYr0qfhGHBJ0dGTaf3aFmE
fWJY4wjCWOEFL+IlFoDZy4Je9xy4GtyCRieY9v+QjDbAYVnPeO/jE/SCLVm+MPvn0Veh/uHvk8or
hz540bRpph2wGQGH+Y0CG5cmUXyXKOlvsNFy71V0nPyT8wtlbSf/idE0ZVzIH/vz14uj3AWKB8LV
KcysqtMpIrfEkXUcJSICICoDXlLUhGxn1T9ttexCc/wZuttrtBIa2sU9GOcN/lEKSJAsn98KqmtC
Fs03jrn5wHgHkQoJREEySR5y2SfnZqBOw7eM1MUCFLEXtREIqZ9fyWOi5+ImGwttmOFXgu36PxAk
LoBERV2tz+/0Y0Z+2AWSI8M+BzZCmksSqhS63GJ+utiNoYnSeeP/ugUv/c6bgz8CNDRme3lQMYBO
Y83hkr0s9cDl08WcS4JrWTrSHdRwbjDH3QXUJtvlEVrqCh4sBrZnDAGM02CjhG7Nk/EZClV8R5zq
j8MRUPN1U7FH7FVX8OVJ7pK6ZMqVyIsUkfOnoPC04Li3TfU2qMgjXbY3IqqrCt+H6m0urq/MJzwT
eAvCUax5RoIDNYHH4lLpZ1Ag8vzInKrD/kmdSM97EhHt7Kuz+JIg9pWmVVaTtbK00vNNeR7rdqra
k7eyHRRPQT3jt9gxebaEqT44nE0x652cWO3g0M8RhjoZRt150Wd2h2HNvWfysYi51IWUaz6DjqW0
AD72Jw7Q/UuyKFJg03v6RMrP9oJwT+e7k+dsRXtio2CVlC0d6l/+wcootcGIyko9v8nQBBf0iDQJ
xZN53vI6wPZCB/vytz2Z9qOdmi93rswxjHIggjhIITh/4jxZB+sB+toIQ2V/Q8pLQoMSeuiwRQq/
AfCl/a9WlTuT5LwA1lIwMexikYBTT7i4Sv1dyKkmFqLU7MwTMYGcFQDwdvnEqawi75frNMEcDa1k
rMhUe279pfmFJYBoXsYzSKjGIzay8pwPrcbFvuq0jgb+1bbzwKN3dIHrV69FjpckTSmA3SirWSbc
1bg25BkNA+PfpvBxRstf9Ba2fbHQoGVedUCTLvDT+tKj+PZtqjyeqX0/3JIhZ7m01gaFykTFvbDp
WZQ3X/7p48NXW5MlLqrXe/wCQ3I3ZPQykP3Vxzhxf6QB5MErhj/fcn7ErPY/iaiF6E8uN8z5x1fI
erf7VnD3d2FmJiH6RX86rPgQZtlxF/flcAhiHw5gG+zciNnmnrv4/LQzAgYSrmN1c57CEVMUn6Zl
V7XP0/SSllrPTp0zOGEtY6sid0fbfHQYuWVeNFeGw7j7aeuT8GoROzvB0rrinUrbhCNIXv+xlrkS
OcyYNE34S1/USZhZFKgpTw3nhPf/nZyra715YgkrQBz5rSqKR+6gh66TFZgxXK/Sra2UWJ0hz7M0
W6PQuKpiquqOZAc3QuvlbCHxSdMdTEF5FH7WlQf2r8bZffdaupqIpsojXfLEhPk5oS/oef2RHzqk
zgOd4DELsfbOjRxeGcXgGZBSoCOSrP3fWrRUxnViR7hmEq/mHrPtboJ+zcu2ThrxDSXN9/ruFQzV
8uVfOITVxbl5AS/BZIsf4kO/qm7qETSZzo3tBOmlhW3x9WlFQn5a6fNtVdgrkGHO4HOEhRwz7B4Y
WAvG/r6L2GtuxJyxSFCF86/kouqQraKIbeKoOsvBbC3CxBUFSzT2zk9XtnnhtNspTr9Evce8hfwv
Y53N92J2O8a7GMtWvT8l/A8Di5W0O/qPqntgoAx0gBbA05wZG1F4jqQiAH805nJxj6u96W8BBHIS
DDQr11M36Vq3ocCk08yWOzqomODbn0l6Cj+UAudXEJ7gnmb4k72JT2Yi6U5E73e8QM1nMLz7iBmr
hsBjEjQGsvf7TO3f6lN6E6DuIlyPTpFiVlEQ75g4L3pWvOMZbDMWUOlNB0loqMOrkgFLqU4ugQZC
PR2kIMZdnTg6+gJagA84F7N6673lUMrfitmjIjsjHeB/R8O7xQyIudDV79SiAsW2Xpj/Fuajsw81
SobpWgRLnVA/UxJUYu7J51lCPla15Kre7dQCSRGDssLqMM5UztQYumzf1wXG0/WOA0/Bv3FqhG88
bNcHBg72FfsfHmOQcbBgE+rDtcaF6uckNB9ws6vUmwWuxBF/8thR88hiCoh4dezuNT8VKWNpqbHY
HDWT2KcjHjc2xchcbwTloeaxwEsj6txjlQRdmdmu8LJ6garjjx89WBHbx8k1bH9MY4HvflBud/PB
pxV9g2y/WsMpeA4AM3CAa9JV7izafxgznmO1bxIJpZ6cmKGxSRiajjb/fFSqBIn4gfOOZsaES4N8
aW8Kc5ooTZYwvvbeJjEGBMa0gz150DQXl7lzFrqlAgkThzblT7vbd2LBxtCTXpUV2/3lBeTeQPHk
Sj14XzhdSjt6QhIDOIvnckHXVPwZl7+XZ2El90GMPGa3l4yp9w5vWcJhNJRSUC3/Hi1vQmxZFLUK
qqj3+g55mTuLx6rOwDumI1qyK5B++4ToHdCQ+KY9grGVuSQHOvSgLnm2oR80r9lveraSlDxy3Vim
ha7XPpxdm78r0qJ6D9c7vnoe50YkFK5R83VWl+jQoyTQLuK4O/dZTAIp1x7jDenV8aQhu/1OzBAc
/gn1RTHovKnVKvkR3UJSH3qnvzQ0O/dKNFZBKzijDYZUzaRzumRe+9Cs1vNaqseTNgr8h/Aj5h6q
AAAYDAV/nvYK1TiFaUFAwSgzEm8gFow3NiQ/YmHML4nHu9mZzXC4pjdOJDkFwKZP3f1a/S2F0khW
7m6S5UVG9TzAbwgcvtAvm7zXweZC2i/Znl+EKil/wp1K7Wa5rN9Y9BsEQsKvTcWiA9KHc6GgVWPG
b8cqWLYNVE8ypmAIK3OAJgwae3/6IwePymLuaomy8vkFT49UJRZb6WxnIvgxx66YNPoa3IUiyVZz
qFoigWL3/7JcKZGuqThfz3LnJoc9omwf1+FakOSdSN0YEBL1ZlBcaAZ+PEb6XWVp60p48lVD7j7z
rUWanD/oJ/ct9HNQo81aUo+A9wnjWBX6MYfGZmgOkbr1H4FaDM6xi6q7nBH9q6FBVmGGVtaZ/hx8
GJX1kgdD6elVpQZ/7fvOTxxlXTuGZIylrsv04DYGc2u3spXaFd1DGG1/JRZUO5qM/2iu0ZrLdCn7
6uNq9V+Y0Bs5V1VQPJLCImiqvQqg0yueEFSJ1kCRznkAuU+wIFp8b7OJTFZ365JmyW5TD1pro/C6
ADWzWfHdgeWI1u6qI4UnhIFicQeTNk3ze60iuFFlFbMFnR4mORbvItvtczUSCp1fuvEfzXXcciKI
Vcr5dTjAbdyKGP6/yOZOAypUv6ZXQ6XtRA7defQo1Tw7jAobxjY8yfmH7cpuEb6U8ahNYVyxMa1V
g6U4HGPKiUaqbLgmwN1ChdLq4qCXgdIw8hHBb5okoD21NbDewQ3ov/vX4NgqhSgm6YUOPJTYkz+N
aW0oGDXzdSBrExnwpkNKiu1Dt518L656ZQW0VmcSC6imlKQrUi8xyDcM0eHKFQ7QYCqCHiZNchSk
MJwTlJ6UcjFyhivnlRTKrhqYtZrF8068QK9j2ufxksy3z/lIv0DyiAeuw8lqaePZI9mBb/KYW+Nt
ZqBOWYyTXJ0Qla/am+OEr6rhai8S6ydnw12ZWFnp197x91ZFlMSZoe0ohn5Fk0Bqljcsf+0OYQP0
xh7PJ64O+QEeaM2gcUjfm5A6uH1sNXjIWFY0Ep+5PUWSZKjnJiN6e5rs/G/ei7+dJIPIV1fNRl1A
mJC6MbZs78PF86DLnqouvUsk7fWTXV9MmHMzq5ummKIDAZcMm/t6n+7J+pK3AgcJeF+4hvfrR44P
cBTfk+wHAkUO2Cn53Cwp7obZ9yLl8MEQC6sYTjhILv1rYm9IN69nzaM++Xxg3tDfUzKWXlCSAurK
ZBcKpvgE5LxxuZapJBN/k+pOCO93+SqWD9w3RfgBMGj6O8lJwqRPR22Ghuv997cgK4y3GoSq+1E4
wBqkvtr1KmMTmpeM8KEm7plD9MNNNU5t6zpVdVzjrOBJbBYjtnNALkJtXEYw0oEv0gZf/oYE2BfY
FNS4AtIYFvga/Gl8ihH5dGFbZJNvzFgWWsNnCW4q5j01Vgbes00EyfYL8bMY7NjFXi19TjbPD4Ud
UT5sWhhPImxZQZsnO6gJTKausZ+w7288dcTrGjUVDynCUfROmq/6Ls3E3ft1DpGb4lUA4DQTnz11
zFUvMyYW1c7r/oe2FF2+8kS8z08hMskWssQ5Lo1WQTqF503Y0A3Btbb4DvjXd6n/5mpkI0NIPU8f
SOoTxm4iJThX2hfHm1AjvUSWSLFnUFRbaviormz1qsD2I4jDPes0/Q0VOQk1/HDQXv5rr724yfxU
6qYMQH9n46xpRdw4T8K6gRbRSDB66aqD3aRuStNNnTA+7YAf/6spAXjKWVwOoLmONw1Y1aiZrQMs
MLEXqxvFOsjIMmKRG3C/dI3cJ89kqTuiuMZqE0nvOQ6af7oA3oxqvsCTLfM7Y7Y0oCMRO8uvkFNu
n2FkcD2Dq7PLPgZsqrb1sqphQ+Wnz8EBpiuEdAU4L75jc7GbNLbfLxhzemHKv9eo652E1VEcPgx9
DkprLyEbZL6KS/sF2Pgv3RIoLb0fD1HoQWtS6WPcgRpgRFINqIgUFu8VOXO2Yt1alRuABqz+a1Jm
VE4dCQjsN3vbQEbTIWFb9ujSrUDlpgNeSDyuVADsHnt3apkZogrYsMfiRYFrwSCfsKuiz+mW0RBd
NkMvGQt7EsBALHDHnxliLGNOboBtSuooaYO6ugaBcIk+u6Olq4btojNJtecheB2ehVJ/BRIMhy1r
wjLbZ89ZLT6DmLTaNqmnRJJqwKBgzVZadQllcyYxPrLYkRi7jcxCewO2GN7+2uHOeDGoavuXHsCP
rWOQfKEb0naHEhhJbQ8S2vyuLblDEJ/v4k2IFNYXyxR+Dgost4CPW1WRy2UWAdQqq96hBhfTVEuk
geFFWDXrTTFVmKGpf3BFtzt6jm/b0Tc5135GUNxJH9eS9oyIFYVYgehsGlvIlO2mggmHPVBcid+H
fDLDwKG9UBr+Fv/ZRB9lKxbFmhEFlibjKJCmhnFzFKXaOQl+M+vYtUMADN5XgJJGmpqW6CBgTqDi
ZOcbpfjGCFBZh8Ay4lT06wcmiZEbHysK+jwH0xPOv3b268WwANPcFICI8+efNCsqIhNsyHlEJ/EN
HXdjuvQhwpnMIZV0dNaKTGnOcWdM6TIBE1k++KtEtokyyvytRi5OJWznMEjzKHfM2ZjzQfQ4xBUz
l+fpwkf3o5OJiRIRViMaYQ1CKRg9mq+vodeqZt860Hb4fVGXao2Qd5V81ns5Q2vF9G9MJ0yxTO+c
7L1IOPiJIJP4WDl4NOJbsAwIeJUzxYrCZzJGlxe2/GJkKKq178sF/toN6dQU6SAvrvykZLowOi7z
3DZ47FrIcqnJ8r8XsDPYsLVeT7HWVCidWMl0jOC3bdg7c+JZ7Qawa1zgRwYCMvgCYpg3IREpO6QU
3HBRZde/0dQZokndBLoDb6GPasaHkmbybSCe1mLyNFzftmc0Eezk80paMHImkG5C+8XPQAN6ssbB
7OutEVGuyIZtdtI2ORWTPeM+k2mmpZyOunZNCiGNNfzjR2YwH3/gkDqiKW8l1Wir7TcszCMeT38M
a3Hqq17tKzQFy1gSmc39Un7fw+nubKvrMsGcjayKtq4CbLc9Q4Z/eQruFRjWTK4Tq2cTL3Zz8mxV
yVQlAD8hMFP44030AaLJNgYVOJkJ7AzJUFm5KRb4f/dhgS4QtXXIsM92ZnCJuR5KfAoEqF/A+dMz
C2ikkNYl/7r0ExygDVGMGjKqLzWtylLamz2p8cTbOP+lKTQR87x/3Q67LKykB9pihfe9AbABfXWh
4aRESs39hMpPr4sEk3k0jtbq4yplGX9WCYzH1n/7oaVwP3bzRQQujIo4F2kP9pO6Is5hChztC+bi
wQSLQNFlhDWi5ZllLu9mWzd3t4SuDi7XZFBfnx8Lxy50GAgPN/ZXxG9oJW+pBbn0IFoIRrT0KAXy
EgC4BZOnby/u7gjv5uM1M5+c1Z9aArd6tHtgc3TOHADmLzfbZCWBHWMuhNG2IIX8mOsd44vKVqKG
no5xSb0PGrK0xrjXYpdUjt2Dld0aLeECgUOGFBBeP+EzFVxKRGkicI18oCU/yGhE92wuHK+fTA+o
cLECSK7mPi7ldjCNL7bzSK+1yMCX1O86P5u6/aszU/XGLWtvwZamQhnDuwxkMdwPIHeoW8kbFydH
32Nm3ccBicsEM2l6u4ztY6NHBypzt7PIbWEh1KIzze9dB5hKA7NsMamVod5u3bUZAtVNcZUsovom
z1ufaO8H070SNpgdkn7e5bNh38aSsIzcZMD26bzQH5VjjJtN+fW1NVkxA3miUoRZDQlt9GLGEb5p
qHXDwlA8BbcPr4vMQO2ClCG7H9XjHAdDAWqZAn54NnXpl5MbzT7GslKyAakiGqjdQzf7JlReXkdn
jfhZ8aQIDxg2wFmvNU1r2AL3urYNNBT0WQbZtRTSFi4IBin61eu1vB3MSGAZOR+ZlehVeNM2NS1I
6Mm1jrkhaAxE62FDHkIMiS5GHHVivrsqTs7zEBNz+AKWp9yCq2tsxmBWFAq4fcr7HVMVjFYWWKBv
scCxWDT16OniJUM68uNAzIZdgGppvbgpT3gWE8bWDjh/FUw/DhsgOSrqe+/ecIaviw40NVB8C+ct
/eutKh3HTb9LI6jvj2vBQzokvpYHzjUpfmcNTvC0AX3bQNkzf59FQcYB+r+E6Q1YgnZ04oasULqB
C7LBikgQhzMQTcLboB4ofOB3crBD9TLS2EB+HnJ4TnNsmTXCWybTjtcWkdRoYYE86OFaNJqBDZYi
2+QrbmR6EcwU5hR93jJJl1Av3BziFApDUS4t7I8Sz1i/CIpavmcUCKv2f9TqLOZPfrrHthnLZzLX
tePmRd9D7KJjFhx8RJ6Dxg/Ogi76thZzWjPmAull973AOuYzgOM/bUhDkzjhyFWgU1zuLPBF6Lya
DvoxcRyY6PUJNkZKTeZAaP8PfgSnYXpDVaKtmfbFMRom7qqGLd/MCzZmPdxl3Zg/80YEU81gnQCU
qbkSPzSQ8sjRrVecKv1pxaWRF2BlP61qS/dMpN395sVvqHQ5JEUDVozyWczsNK4L+OJBJAT3naXK
CIuJZQUEa0W6VwSLxXl2zQ1g2RRYVFImSU2DIb0LC9su9I0W+PZdbb0Y51AGUvEuMajjZaO3bU6y
xwYzR9xK8AHlGz8xwxMnVTRndahxjqhcjgD9K7WOQNmaNmz1pX7QQ5t40+f0+o4FpRsop+ZS0C7N
/HGPtNBd3ed8MWfHAPszZ6kZf8BEgm5fVikx2dX7qTKOnuq+YLoPnMR6fA0QlaC7IwUUhjXpj1rf
y4IWMaZqUVKsPKwYlYx29nyaRt23jNjq2v526JCE3mqQnfKicDhrD2S3ZPrJ0IgMOQxFjRgLhok5
TlQRd/RPgR1pPewLixfMpLhHNHULOUIzE3RXvxSGBbGHTZ5fCsCJQhuKWwlPOYiKi8I+JJj7q8UE
qWVS2nXjsbZ/SnwRNwm2vEzEeSCrP9EVSqUfOvv5j2u0tgstkv4Lr3pCrj019C75OlMOa10QrDQy
qfkHy0kvt1cXdcdUM7q4tixrz+esdjLtZo4AfSQuRCYXHn/lcYvMLi52yZl4QXuSCaqRKqGCndVR
CJijd4zzxRpEbbhIp3uBrJ0i0tRBB0xcZDyDWv84Nh7NBIuJ8jAjomXwT1H1+K3dXZ2zWZQiB/9P
1+x9UvWvWRokXJMTvD6Jcn8e8LC+7X+8R859jK5afveGxuMLyakfuuyBOsngwhaA9NNh9qcjNhrA
nOcqAJG+NbyfLwVc/bZfDG/ghcU8kxROB+SM3cqlAKN+89zfYWOJVvACWaSjG89FQgDmTXRjX9lF
MYqiOB8v+weOEhXyEJRVEEXOuFbjXIp8s36U6sySXhN6Ye0UgJ2EZosAXsj4DJ1nuo60f6nYuoBK
p2WZNs/1D2iwJsuYfyCwLP1cvh2al2aeoWkIAmT7ks4JgOUDeYyeTcVX4KT/6ICaJoQPcy1QG+uD
oapHmsmAhj9+SJ3mOyFunbQBU7mD/rLtUmDf9ANWs36qzEAjg3mW6zKQ23KCj95eRADIAlozeZyB
j9QGdrprKYoqj3R86hZMkE/oPDTMpuBO+qPMNZftYTwS9XuFWmy7xWVqEa+DEjpHzg48jaIQcOF8
3GG6R1c+FDHUl2SP6dl7X9MO1FqHJQ2J6Z2dJ29tZMAw4z6DWoAiHvBx3O3RDyyyl0t9j1fwb+F9
yMFzvxnK1em9At1rCednPqnFNvYFIkwcjyOFiGsKTljBdJTPIDMV3ZgrPsQvn+phihdz4L2ecI4c
Zk3DQCXcnK+NP6q60GrmFr4IxWm8kZudy+1BtUkVN5e7xrmgjAHeNqM6iOJpxFa48CEcuVxS9MLZ
RteGiPkr5xqMCWLTU9v0Uz/pd10WmYGksG2OlSbkENcODq5JDZyXXwMmBPcwD9LGPwQ/8xWyZOQd
Hds0Dfs7sxspz3CIP/GP2dnuWz4hzs3M7Psk787mIu8jrtUxJlC4USkXhYxSQg2n8pmfUfFZUKkw
PBcVJx9EcW1EzbLmatoMPO4ke7Fv5cZnNQrmWZQzGTIp/Kd/Xxnz9I9x/LjIY43+O1jl9MzPXI1d
MgmtDSitv+UQTzGq/6AvFz40ESFJUHSykWQRgpCPERVFH+dNvtnCN7yHqYZbwwcZ6kYGBT83kCU9
yOsHC9SXlOuMsDbe8zWBzrg4GPtxDlgPNj8SlfP9Wz9BK1N8lVXlQqo0024jjlRTJeEA45sfERoZ
ZOMwPPN55/B+RXX110RuV9NQWoPcDq7rnWP99MbRN6trtITSu6CUVTd+8aElxjNIpxIiNT0Rti3T
66RzGvpVT1YxVcAN/XTf/WRyFulV06L5bxktAk7zI0I1oMqd7/1LfB2ArcHoU8G2XUmAtHflmNay
30pYetBshCixsmyvhyx4JB3Rlz8dfatZDl1mY5bld90iCXgVPnrpZ1C5jMhfFzC/7LmivhbnMGVi
bJ/3RatJvvFWNVwbPfv5R26PKGxNX8+62aWewRaAuuQ4q0HfZtwFPGxXICCIE1sHR4u7akCH4N2U
XViVg0roHIBoeokdEhX+BScet3uRSoXWNhLT5fGXWmhPfuZ5sb84jORSPIrABBqcWZhauBokM4lI
6IcqiikAlUYCvszpWUQ7yb3i0XMr6MQ7/JpZFEGoKoVfo/54Zm2GdBLjOzjrWIKJErguu3uJkJRc
3NDbRZIajtam4AG9tr555bsApPdPyns14jS+8Ppn12t6UMQYLAWc1xzVz/s3nh1qTz83rg7p5yFv
gqNeGjG6PoIuQclgp9gSFl8jbjglTLURpeDLgjiZyorDQX3qOawU8gvl2LEUiN1v+RCAXj2nrR0T
HOvqwmwvScO7PZEDPhb/N6RSeWBMbD/z5LRZSOf3ZSPbEkLEVnQR9iDt6x1S9bbYLwH1t+oPRcNk
0D3WCFlaqsVnmqqeiC+u8I0NdLAXuljQQFx30HbZC1zZy5Hmg7IECtbFFy42G6uZ1G5ORZeGtrqD
AhZiqoTFtuBlvuMDiCcQJ+3ozObl766er3WsG5pyQ/wuulZ2MIfWg6c2yC1xu/cYpzRs3opepuKj
raWWUf2fRPIajDiTfENHnUgwRsGc9YdmCjXN6uW7g5IiLOhm472caEyCg92FcLwcmzXYh8aXzizl
vjQgdncBT7MPJVbhrlmd75rlG+tZu1A0TwMoiJeSimNlnN3HL61/eTjtZeqSwQPNj0ndRKt+yu9C
UB+gRR2GoSSF5f5JXvbqcyGsw1YjMI11XxF3zAMGp8gfRnr/vH0eBAU3u2as8S3aaLlNavMW/sjg
l9WhTqf7wy12orue84umAvSdt9LdyYwViXB6leguA14IASlABDmh15mfMgWw8bXMjb7ZAfEhhVm8
nHVUSNdstGgdgv9b9vm2hqzvLb5bifNqfUI4dvyZphNKceZo1YDqDLCtLSBUWWrnhC2g20ee/hnO
RwzR6E2C+8eooMe7f2heQmgXTtd2KZtVGl18GofGA2AQEAkohE4b0xIdVN30Rws3VKhtkNwY9nDn
+vctmSWx60eiDBrlWOekeSDRdO41vFqO5eGc4I6r1/ekWjOhMV83DEIdkDCjWJ7FpQvoCjw4bM4j
+Qmmtzt/oINN3pkXqRiC4uearjqyilEOXzBYM4kHeHscOItpZgPAmUd+1rSSjfKIQb6u2LIS41lo
pADw2EeOmtYy1pioxQ7ubzr4qTbvNBfHyyo26pbokVjSSXyA6zT2SlMUZBTXB/kvGNyBV/9G6nZR
od6C5p0TXT+emboEy3SBgw4EGBxTrd3LokrUwJSH44hxpFtTmICBdrZgF9TmKcE/tqtMp4phwtQj
ql3mLYmTJTkbKzRpJDBW+YKq4WNjoTI3+wHE37feiQrPpJbwVC/KGi8qoa3bz0B7NLkGLwroj5od
u1LjeZ8mjkWhYm5cfM6rqm+lJWc5Ep2s4Yzxf1xL5IzcEx6V7qLSHZ312xAOZZ3zLzwAlh/Lgaw8
ojGQYMtVz9ulXsn9Mp0LNbg1TiT3ULaEIIIs0sCBCAwZTGDJrzMqIJuvYgUsVy4/yahbxvEt/Bjx
uy4APkUeF4mmdo11Fj49kQimXebG4UNMldUi1+t2KkVKRIPlLLZNTvsrCYtZpxtCjak0d/anHQ6z
x282GIWGx8kL5ZV4XA503tJ1fX8Qw8VdaSRg/HT3l7eZFGJeezWYQ3kMBudvgbaLs4JP5er8DM0I
KWWowERpWDsrUnOAYK5KORCDqH9KaD05Ne8hJ1BwjLKItSj2Ntb7/3tfv3IAc/OTU98GeGBlmz4v
eItzNem//MZVZNWuYqDcfkqPx3WQYvbjO2odY7sSF6MirlD5Yiw3lnYVzYlWblR0HwCAVXHYtt+4
f2IaGdFJ9OI4imBlXbNHVFWr39o1jNUirOQF1pCTRBbeAjDPuamC6aRPMYgnLES2ArPf8JDIdDhp
toI5gzM3FeeVG2Bn78Y/14ATPwN5GlqxfqQvh16Rno1t3ng/E+WdoeqqvUL02SOC9cUTAib/JmU0
32tlrd6IhxXze5v0b4U0Ey22B3JpPud1mhu99zOtcQz+P44MyURRyqRCaify16ufmaoprxx5j3wG
8WVhx1ji9r2uAoGlZKHEVPMwdH/sTScFLATVKIrRhTxy1ikGCxNiG/JPqSKi+liiDZZeMd+XHyn6
UjG2uzTIEzxwDhKeqpzmad13Qyr2j44mQiv0FG/FU6Xrq9ZucaVCKfPlqNr4XhHLMV8VnyRUszmr
f/IZEKys8Jdxj6yWsptf6pvcEKTExxqHwXk73n7UZQBbmHLEFYUnWA31YmotW6oKe+WpFbUlwDpg
F6XikvObXErUvH0I/x4FOPYAmG6fSaDM1mVc5Di2vKKsqAh4kfNY5XolTx+6LHZ4rUsj2XuWD2Tx
0TyGrEF/USBgO/MfYaPToO4P8SCTfQPsm3ETj7drj4PkFrDnarMJS9xT3mUMSIeBoMgde4+5QFae
YRVNXxiBhjVO7qo+tz1Mvq/x9lW770E//+NvIs3b+YoQ9gKwK5UbVHya/dj53Vr5wiIzsP5B262K
XqhH9O0KkzLj5Ds2zYTTayJkwwjLmbyJlNobK5eEGpKlSzCXSjzLFn9S7YX0ZOvetAPpQ1JB0eTv
qmM2g1u+bPP1jw+qEt2ozb0YO1VbErBN5RPYK+5H5ke5pbWUfSzIsX5PGZGdIZaIj7lEvLgxzThc
u67NSWmEE4ARLjz0wfgKPB+cppj4kv6Awxhf7LJbaYgHjNYKwYh8G+pLuIjpTzzG6TP9BUAJp0bH
v5v8XijXfHUAA6GfoFr6nKa4y6LgL+i6M9d3SkwMH1UpOn0eOedLTBe4eYo3GztylGsHYQX3Sl+y
4ZXpZ0H0qjVdp5WkaqlSW8mTkcdhgzSme4/m82Z+FnhCBa1CMIBme2q9T5mFmKq1HQvNi+/SRG+w
3ceoC4ZhcgDtzIecgbRvonfFa6C8q3L6bo+6bocx3FU4YqERmCOx0gNDdebUYvZsNjCHv8n3phAr
n0mvXdBhh04+5g17LvFaCwCIaOfXHRJXUOqhlk1tzOyaHRzJ1SGH0jZLkzGspPDyIaDV5f+gjAdv
UFbBtE3gaq1yuvQyIbpk8C5mSfrk9HcxWwYCqKB95zCSW8SgWmYqWmCBSeQuX/6jyAxrS1Enxsgz
U5HZNwkf8vBfwi+OZ0KoT90azY4TT3587WbRCntb2KVjJDn0YTy/oYySOFqdzj6MbyoP+zVvTp7S
bdbD+7/ETMAQEFk2thWHC+i3pqFKCIH3DnfxO84lZwCJ8ilkVBlHadBsI7XtnhLfwRNiFggyQ6rO
VcBtEVGEYn11EZqnKp0taUscivJEXoPtdLoMuN9vASRv3nr4am2J1NhifLWrsULJwyqm56cptccQ
RCRJHg/ua7zAMvRWrfzWl5/VFoW8p1Zxe3GbdeznGxH2StxzQ+d4ffeIFHGFiHpOdGQMqlTeaejn
5Eva7qXYV3FlmWfkbNeroBPYCyVP0zALZ+mia5+cEf0wgxgrx9Pn64lHd++IxT9PZMG2N9pD49W4
BWNcbHPEu5MOK4zBnLSG0/2qC+0mfsysGm8PUUYCpXd2tFJlyKond6WpJYKtrr9/QpB3KoPSP2eR
OF49+SUpyU8OqyqTl8Du89BaUGZA1rbtWwnzRhel/Nkz5+NJPa1OMRhulxbSIUPRg3Yt4diK9mrj
ts+LGfIMUUU28fduvZBzsL3pEqo/VsfiCXcPZ1Gt+tNDAgFJYy5sMJRvH7s0Mc+srbePZlDTfo47
dm/axSWoBHnHhhLxMCLBroASkWLIw8QSPkiqdWbcsFpMW3R8ALAcu0kUT2fqkDJg5QiNvLRNeXsn
7IiZAY+gW+qeZRY4RXZMlQCW19M2ibiaNw8HdaJP+p7k5M6+afx4X2OQsio/VVc+qB7hnB+DiZLg
D1e8eMQqAZ1u6LFz4yvTdYO/59Te7/8CHJ+K47X+57QSbPfNIlyr29E1FyEN1ZMMtv68bxuWJtHD
9USYbHbzTwybekxxx9zVxQd8jCpwhWW1J343Tir7SEWtbLByChcYJnUgkiRpFqW/7tUFHihBVFPo
fDLFI0vVGtBMfBxNlff7zaQtaUkQlJhKp4UWLb7+PdrFVEBohDML/LhWItElavBFmWjHRSty5Q6R
BZJnM+v7eeS5ngP55PQqlRZ2bZPoxSUQOuoE5BrxiXHeGizc2Pj3R/R3Ilq3zHOWxakx8d3FO8NO
p+an389dLZMQ5a+Ds4l5Pi1v0BuGLmA5UaFnPfwGb9KidLQMNOvxF8bAMon1NC67fJoBHp4Hm1zU
odlDe0h2ux/Nq/NyjStfeQ51WvELKIImU1NTkuB0IrDw5GNau7W6VY8bqf4fI/a3kW4US1VuO/4r
IX62XxBVnWsnSB4fZHXBxRn4jvVK4oP8DNZ2IPMrIyUycUarnRBbytHpsbA8I6LZCzbjO+CxpOqg
0/WnIW1LjU2sZxjNfV13Zlee64nyRhCTA9xS/B+GQEZDjR2hhw0nP7FRA6BXoCoSYzeoGGcRKVKU
Ie05ETDuTmSgZuMNQ0AxU37JJe4JpTzE2ZXlOz1aY54OB/+JG5OD2CEuI+twpJtl4xLSojWhiy1f
keaj3QKGccg1E/CKpVwIOhUAgNBSmW68ZIH6+JzEDRhSSdK3Sn2E6hT6DKWhgXrfm3h1xILvzXHU
iCJ3HK3JJ8XAaZ2E0hplcvvSJjmwGQMTNTnqGu7u1nbGdD56x5fOki+NYEldkKvdQn5VJsbgfG8I
8uxeOh9dlKwL+8X2KprxIsBlKc2GJMyLtZtxzk/uukJOso4Iqb80mh/5kfjPC+BHkNWTwrUksqIC
ebd9Ju/chR0tNlTL0WJZdUS+qeI5iYSoXwzE9YrbMH8zqU1B41IKSC1ZX5vC40cNzu7hJDnrb3sq
sHMztOd4TESxbinSXBUVJrRtMEDBNNSBGxGGKtBH8Hc51LfCC6fTevA62D5N3OAmsmRqotwboFTz
luyJA9jR4WATEMu+Lc1XqJlaJbxxmnueJDe5NzstIxRjiKTCjW+AFqMbTQ0TczHJ0AUmIF7tVSwP
BCXz0oSjevWptd2UrKO33tD0qvzIz0diUwt9IXF4KUGx4gXcGRK2+U3gKpoSbhUwyz8WLxPyR69n
4lAb3guZHUHC15hijo6sBjrvbemwc2jtcCtJmmYHrh3XAfYWPN7fXz8LBlRElL5gs314XCcxNVCy
Wmueyc3kiOo8FKkpoR76nlsJgcH/tsB2cCxAz0cAbmQUIt9XfpqGHnPRrd++Ee+fH2neKCzb+iUC
qFzOUcxgwXDUEVk7hrEQE0okzzrtEN85zwAKFuD/I4bRN9N9wA9wTekMM+gurierG6vwHjnuM0Y2
Pw+2F2yx8f/2LDjr2D94vMdA/cz0gn1wJOIVP4p7vFoIoF2NOGHeqzPaS2LqRRfu4qxBWWTZwe9a
Xt2n4n5tKD9W6dyJoxYy6glpv5TqhO8a/tFCgnBtEbxYmLOf1X6OZCKV3tQ/f3BPk7LCKYaMqwov
6+L7Xt+3KVQ86KtH3QfSgR4QFV/SiXTMaMUCOex8/3W1ryvj0J0CHyxZ2/jNzcDansA4u/VEChPK
yfs0UUoKWhqjA0U0HelF+RWC7LQCDfloY0fEZpLki4MnHcihmW4Jkh049gKHIrhUJclFDEAUlpFG
A0h0uQyOO4QeUqgKn0NVy3cpO1XXeDjaI5d4cQX8ut5j6tFkbiJI4/rQ/yeGGXSP93IoMAiLvm+6
3Mh5U55H3jeQK/m+rw1Xl3i9jsue8cP5xhkwJ+UTc/tIO20yhWNj5NtJYZrah0+be+D5I7T/E1xp
wJ77N66mDK6tjY7c3P/oPPCuSBg8onv8LiS3NSBU0Z9Pa9t4EnklP46eimfUNDHwL8ipGJ6lyuGb
UaW1k9H5qoNtRp6JsMavk1Vvdm8e/cnvHkwb0wUgaCb0ohzPeDLFjETTSEy1xkagLsegIV2LKKuN
cbcynOpyG/ZCJcdaqi2tBM+gG+Nc+3esLTUOpfUGpC54vOWQ4QHEk+pYNXxDMkCtSWQVDTj8epZz
Qy5fIx/V/6tZpZSFjDrZw+Q2JGfXkggzJqoQiQbdqFhCHM5Klyix8RJkxdbwZSlaoLNrwsXQdv6D
Uz62AdoCJ1DmfovD0qQu8gfXdwbAyeO8eAQvCj3SyJTpJYbdA2aUxtlkvqD58uAONtaaHzLHR1+4
pb7m/SYIsK1l3aFNPaXJo9e9XTl/P60/dEpOV5GIDbCIFlm2lY1mnLiqlYXXFNlux7bEQlRUu0jc
2jqgUvGonWuDwDUTgTq/XiDY0gUbERF5+6xiHQfhi8nk9u3UF/R99w06B12QNnvDdjlVRJVnc13D
C1LK7ESVaZY8i/EN7JMZZ0yMe2z3GQV/7hUQixfFhWQVSwWOwp6nLdeH3jhww5F9aUYOmYprLKMc
mA5IJrbWnEdeBWGwJOrF2PbmZ1mbEFFM7W4+OCBR3Ty9815j5kQzcYZf3v/JGQOjFDl+9LrdJQJe
J1JEWjuPrQybD2EXK77iHqGwPw/qErDKnm4514hAofuBnvLJlk6ihhwlgBszR37tvKqtFTO3Q8sk
AE59szXyddxxdGQWLFGGR2KTUUO61ebpKvCIFbX0tiKyWtkSLUV+eQ4bII4JBTkRlHzJN89kCx9f
dqtHJS7i40j7OQKqRM6zqCJLeIr9p7YlH1EByVUc3iYidudxlkk1hkcKc2/bRL2nMkNldZhFlcdm
Dy5/OMfELbTFrYG7qf3ovSK+fnKcI6kebyv81kUpTKFpjGUqqbtSUIabxebtA/hI5JghrzjNfcjx
ML3CKwsOYnB0AbwURzQ1P1o4O5lBgy2DtmD/2UH9Lt8UElJcOr5VHmruIs3enKpvT2SlJRNjNFTr
gAlvnS+wRRnktMKWytcgk4zn35/ImV+TTBQp3JPpDIxc0AkWguGVEDMwMsHqZuEtCk/KuSEAM204
xaZ1UlbFxe0PpnfdxUiPZHS6B3y+uwlOOgwNAhye32y+0zEFgdo91r/3UPQNxwy08bXFcJw16o/p
jjgiTVYZ9krunGdqaQmOby+CD4Ga9NeTy7H46wHfdUsf9Y0SiBv5Jw4DsAXaXqPufvrXoNsj5GQ4
/INy6sLgTpwo5G1baA1E36Tn2inI7CuG4T7u/mMnLpxUTFUDb/ot4bqaE/S3mLOPl9MPDyTQlrd0
JK0GUZfAcJ7UbmT8y5RxfzB9UfjnqiKgwtPCpjnjgrpK8kqg24jxQL7waaQBtop9i7KsZnroqrTH
KVt5C8LOBSQPi4/cYfh09ZK5nrLPNLAS377wkarUz0tpGkYloDrn2uurXSqs0SJ+/WBUR1o7at/D
ccxvEq3mD5V+4T5dLF/PBuuoVwb4fYlCZbxg6xDkXDy6WBcVFU/x+DkeseFakTro5lfSQwyvMS7E
QYRJ+n2R2hBtioqI5QyN+X13lCf6+F6+Y9tymcs/V0yNZ9zyAdg+q+PPYgi09ER+PiM0p9Y+IVTa
YO6MedCVzWLrKXOYoMBnl1O+BJcziVH/dcUa+fKNFfSGdqfqps0098XM3ge2thmF7QNqSpxvz2Vj
KtOtMUuDgWKYMOf+FwxQzvI+H/QDitlxDShUaRy9mDDbFzTLv4xzYznpb7Owa7z8yXuIPJijSwlW
V2VMT4SssMlwPn5GVf4+fjUBPh3T3W/0kpnAk7l213pMDLRbCGKEmm3isLv/ooAkt28rSu11T353
5g9O3tVhP9aDv0Q2cWCUP1eNopVFZD03/YcH7a0vu0yNM+n8TBe6ItJ9RR6v4p+SVWGsgKr3hik1
cnn09SMm0/HBsqS1FX01peG9QQ6PWuZmlsaop+hXP0AngmKQaErqsyAosYqkuqkQS39NZOrXypkU
taWSl+LkAyewuuJ9BsqbTW7ehL18xd+/7SiulvHYeppT9VwNPFD5K7uKnB4aiiM717Dwa8P69Rtj
uaUVKu60zyg4+InHl4ezQLxqkb4EOJf6+TET2I9tKKXnc1ZiMcD11dRX/6DyZM7nsginBplZIg9T
EIfIpMT7wf/cCB9vOX3NJ1E7DEQWrF8cwZpT6OKqXfjkeeIZgq5Bzvh1LdOtwkvkgroJu/1yXNx8
kjcwAiyGSG1dOWL8i8Fo8mfc9RqEJMcSraQl4KZCKN0hrWir9ZzPX/JlNycIZu8yzyq3xFSydfHl
3LMXtXsO4LAZFjoEGcyBJeG1I7xBvom+Mr5AF/TtWw65u1H0DpFFZxZhXjTGJ7wJGE7WtmQluntq
Ylytdnk9iiuJW3mUZO5c0ko40ghbnkwH63TFLjOid4HCaqrpeJI0/SBbwI+sVTk0PZYWY0dmdS5c
8a+1y0wlbj0BcMLpu7r7aDGvE5pDHFSxkNOoc2eDrje54CteJcGCC3kpXdkeizj2TwiqIVrx3nve
YEU/DZsSJzzt50n9Mi/avgIDXqBraMjTb9Do0xprzzSFd2nHxgYzcQsHkjgJ0J7/MdHrwdf/1YW/
TmpRsX7TDtl5/Rie6A1nKc1H1WrKvl3fhW6W4GLYIS1lhcBvGAP3ZBLmnENOQ2SvkKuPyUndiq+V
Bd4Jox6sUdinY8QzO5sGykNE3mG1Bz3g+rlanjobfmS1+dZa7k2kyg17xogW/FSM3BCK35UoU6wJ
N02u0QgZAm3khkDeX22XeEcXg0xlEULgcwM5OhMRZbo++FRAWASBhOi2BF/zX3vrhasQKAsBsSoK
UAY24wUbJx6R/Ec+jH7sWKRqrUuQvBcmZoXs1abestIZlF7bKg15rs9xJA7OgQHGDnqqm6L9kleg
Hl5Pbt0ZqAWx5JUNMJWM6c0MD0LGCUvAA5TOGt8GJtL1xOe6zLcwgSBwJsbqrffAI5VReQXLLuPX
xaOcpPNRUHLYLK2jh9GQCnyAjD6Jmb5dyrMncdCorx/XPHJga8vTDLCIqG4DtsR05wPWCM4lfmlr
E4LIGfMyjXqoHxTXtqE0VvRWWrp4UJB6BvNIvJWPnI7qplHEEQSDJtlLD6YhU3BTts07Du0wDU8y
CRIEBgvbz62+wCzWEcTCnbAAFYMKCWuJK9pVwNQzDPVpIZ9kSFGYvSEAAP8Tx7Of73xf+pMZ5RJB
tqnL00WyBvs+REetBSOPxhgM/C2U31kRe/1MlX5sLpKPKxR+iUVUuB8328f7yh77370hhGSnnIoB
ekiR7GeebcGtpi6WCw5tO0aUcM0yNpmnRaMEduEC6VV3oXFxrcW6/gQ3FKdTG5SFWgON8iVl4+4t
qRbbifhDvuv1vU1VudwOgMRNjnnqNgV6GtVhyt6+pLKKljBAn6YpNWRiDd3feMxEPpgVM9EiMfQp
5/jnWKgQo1kWULEMev1xAq2jVkO2SxbIoaw3kHFv5G/lSq8sTyATrvwH2kCezh6NE6U1WE1u6CRx
vZTMHDUqUXcgc+BsOS+a0Z8Wk+vqyVDbo/zTGRS2rrErPo7OQyzwhF0hyRAFSxOInKm+C49KPTKz
c4PZaabaTrW35crzKCXIpdPnXDI+kZY1Z2dzyIc5gkjAv++40fEHJMmaHiilN8hseCcqOE+LHgiK
DShBw6zJuJD59D8RRGcxLQQZqyQ/L5PSUSHuG9/T46w7ntHQUF2VsmyljkZCiImiT+jfQYSdVveP
meVc1tcVsYsZqMeOSouk6ejUotNFu1mTEUzZm3l+M/lyouBOjVGb8t9vtglXAg6iWMIJOKv+RrxX
xeofMdGqQLGN80FmXALonaxiEMXmOIiQuQ5RuwkmlWY1IRoMlV28KSamauidHXUqfaMcrUTOlKKD
tfcfW+0cTCK6k0Koz8Pi7xVAyQOFzUgVany2JsBkRbcP4LPFYl31q2Zm+fLv/4SdgquASuSSf9I1
S5z8pqfW/e/vMljkMzFBVFLPHR7hSlLS2kzOvC1AGOwJm4PIluubJI/zOix3d/ZQmeTer2CkHO0v
rW5CbT9BOywAVDU1YXCgGO1xNY6wsIlwQQTuKpvZlrQ/Igu791BjmHGCVFtFbfz1w2LZ+7+bqziI
5ObwMimpVbBONBkvEThhYbCI1/PFOvj/TOauOooZEOHRxipJ1sLZGPpUpoUSzmhuhL18q4EX8RR3
4BWWWGxbsJGjw5/3TpsSs0waGFolt6mHXzAnPCKrov62wM7syWSqTExRq/S8lNCLQ6K6FQNJSGvr
0tXv1Tq6xV10b/uXmy8Roohi1i4MEXXnNKESDp6NyrxJUTwtXOX7eWYQ5Dp/xGpg87QSHvVBNQt3
6JEzhwxRNqTvH2mKEl18lPtMREF9oWruMhDZMhfhZADUfVoxeMp1yCsqauEKGFIHRL+FZgpRdRj8
bmQ+0HGs/qoYk/Fz46x73XUf4yqJiNQwg/1xfn/Mn+5l5xZl+7KtQZEUS853w4W5eyRuLRXFrGFW
Poour6hzhFFcqe+uOnrACWpxxitIISOK4WMN+ajhAe7QUjUxtBhLWd4RwbCjaS9mTvJxOjriD6RA
ML4SQEXywlhOZc+lKRBkk2/Q+7ZiJIaEfqcKHjG/p6pAOb5cGnMWGj2PzaDyR5Sz60DcQfYOkKXC
G1sH9V24PpEGY2X0uqhXnvE7pVRPOoxzfZM4TBXTGfDTUEh0kyf6z83T3TgnUbGvDzCYFrJikOXd
NsJZ7StoXJLrOXQY9Tkz5aOt5/0B9nn808U4ebT8RvsPA0OWleqpJW6Ybry4S1axz7wDw+zYwSEB
vTLKg4pAKxXDNiW19zXKUKqdsnFyVczxc9UkIzlQLzU38cHgInn/DE2VDXYMDxYBR/CRfHly6etN
Li8nNm9KiqQ2q5rDdvcT5YS3+ImRJ6uO8LKogIPGnVqnrZC9wRQyMJ+SuPiMy3I+2M71eV6gj4z3
XL6dKpU3SzVl9Jx02eBxqDKQtMN4tE0GAlB2iTd1BYk+vTJH7Ml3/46Ly2+C6ij5LgV6e/YFHjjm
P+uxd4DfydzcSZVFVPMJFGAnFBgfxnUGuJJ5vjVc90WgVW8vW4mzdCjV2lA0kgQ1Ey1cG6RcNPP4
brp+1IfLOVEoXp6n/30s9qcEcRKP8WXgarpgUHazsSsTWVuWlCXh0NjZL1mGjplWONOZ0tG87Xu6
WyE7WeYgHNZNw70u3z0WEs4IVBv3ih4xTiotubLOOpyg4A56dnN+YDdqI/8HRTamai/u5NWQi2Ol
FwKQVvMd15qO/3b5LgOcNtJ508+XRgMuPyupLcRbc6P7hYTwfAwnTF43FwKny55RPSpG8qmx8APp
oRguozdFj0P7e/eyGlsRTq4oVGgYJGt4ia+U69hvdwbd1I5aZQMnjoSE9XJw7uFCfUlSfwPGCfCP
4UkroGnO1tJT2+EKDdqw4Yxxv1zCSNJf/f4gA1HCy585F12jjDREtzRcJ25/KcQE0fE+GgoKeNRd
gTK0tY75jvfZwUnFq90RPxuISA/pJiXfSFnSgpGzFOTtkSdFhsahHrBmwM5e1wx3o6ZyKERyrC8j
vKsQxqbimTs7F5Z7vwgm+xJVtzkgrC2GPJLJwu/t2boRRAOQeQ1hQDNM40RFoGKvySz+AwNp3o4v
ZGgIDoyNtMQXro3wlRh6xs3DuMEd2TzNaLUyEGd+VbuR64cXE2cFBamYt7efOw86WK374ppXTL76
ijxMXa4nZ2YJH4DJ0NjR0QI6Q5WE532Q4rjeOlP3HsDpJBhH7qYZb1/oAmKGpGZqd6xZIUIpc8Ji
wAKzqyLsYRx1e6pbAUKPrjLlsc55MDKCe2RosxVd5K6ZPZRzxSpgo8cEldBQELlhsggidqnlD7zj
tGSqEL5goHsZ2HNyFYKD1rekxG2gGq0vDs3h47dHjbt6qJ38Zz/Dz2SiSvtUCya+jvdr/91rupPv
sDyzItpPUNGODQqtgpD66p0cRpFblg4xjVFbzUjgCj3zR1DA2JmdOtTRUwdLpxdby93V7YaIEf4m
ZrkWNlj96o9DYmwvsGyrb3FRb0Wcv9lKGAg5QkUBQ/4lUb6WsP/62tncP9I/8koV7wNzQMig2k7i
6lGJDWLAhkBQl8mGe+F3rYWoLBUWfpwlMQKE2TOozPvsGa95Qemj9JuvBdfBEvExn4tLbPl/3isK
N+Os5kQxsB+BOlzD3BMtn7GgzDzbu86dzYNAZ3DNgZde15n4Q82tLC0YCKJm1WWkUvx3bdz8sT7X
3cLeCbvhfJnxYe8pAJoBth4u3lmXSisbA0P20R6fFQmKz2183EUvYbi6TlUP+QNAxaqb9K8bj+Zk
q7eKf297wLZoErhFNaV2d0zmND6RJg1XE511mcS6ugRdKRFFWukYv/Mi0VazgsU6ea2l46qKSuvC
J80fJIsalJkPAlERkt7MIDumTRMp7rX9TeYNB866FbgVUGH4DFL9A9EuJ8UInUOyYDYQY1cc7qDo
tY0MMd7S+ry8RBaz+pvvWCC5yzoLYaAX1k1XAPsrF68lTNJZdydFWf3vgAisUgxHe4P3waWeN7ap
POJCg3maVEojsXolPJBABPB1h4Mi7qYywLoYThIrBWRyzZcJz4cGtWbHk6JmSQSgANR7uaT2addU
ddZkXE6RSyWVFG62mRdJXWCn5mgYpEapWeDUFFG1msL1q0noYOk8oLXO+0hESXCdctZvDjAFVdUx
lLaUzJrMD5fJPrSdn1DzjdfqrLSgaw9TlkhAxiXZZQsFPVkB8dlMXMB6Y36wrepFvZkZcPwbTzpJ
eh4ww8zQYmp1OHO1azJmLaXLCLS9qc3lod7ZxhJ1J+QZHFiSSbeiHI/WfLGNy24a0QZAdmjy4dwn
9JUYpIEBy3HW4AVe9Ra70Vy49mtGTGnpQZikpJWaziAX3B9QkeMflfEHAvAbXDirix0ZVoG5AyzB
dmcnHh5nJbVrB06uNw9cp+e+zeA3h4DdRoMkAXtwI6VRFuMmTKti3JPs4WLObKCvIWI9uJwSaXjD
ULYCNrovlJNu6BDhMH6eq+NZFKdu23lOd/3CUXKoVAsNSZYOYc2rhu5lQVfYnA9IYg+rqLiyG97D
wMTO8lJKDvSImQsb4x/9eGStXh5LG8GXsNfiVawwM3+NPqpmmYADZXle082jpXG81E+j+ZORy4Yj
4z3VYxoEX4iMRKjO30Ag+MXTVXInfmrk1vg/BhlepAmuf74bN3KS/mVnmZhj4QvrztwyQ4Ma4JK+
78YHtueKe7FjOF2aDr72rAHVU2chHiItdqTITlvDQjjPeDsZFcNS3zfh2zG1X8XaqnVuCOTlILcV
E703+VAgGg44bL+s9PJcuQWMyfPX5mfIMpVJUGVMmFjwja1upMh1GX7I+Q7AbrAsiq8fqCw5Kbws
JcSRwcJ1SL9Q0i1Bejmatez7beHCmTeMSsqrz0xyB67Se7KoKN0hAwz4iAm+hgp+YbjX8m6PG839
AS4o8tffNro0XRas4OfXZF1IIPSIgDx6sNFNWroz5J6HVaxDf8Ggc+3JCZZVEJT5Ntp4apUB6tnn
5HyhhysFptO+fe1NHhtyFkiC1/Ps6xoZixifNsy0V9g6uhM6Gpx6uTJLpfJIIxFKtjCSk2UWqt27
OQ3Q8uD3fisL+q287zPxh2q6LxZh+pzT+af+0NHFmLW6cL2dm3+Gpo/S21v3F4HM+11oTRilmDwP
6g0HTkEvxGOBFA7TLXkhfFoY3+WJpl1reOS1LVoGMJYl9K8XITq79NRKBlGo8haKzyBUEz/b/8+X
QEnwnrs5+wM8D5MLwe3oDZbyJ73TNhVWysG7+/21HJ6ed5uabcxbHX6bxkQt9e0vIKtoT+IhSBWA
dyB88FQ4Yc55zJUxNdB0Zhyvr+SVakmsDI4s7T3O2k6hisUIN0Bzdn2cTJwXP6JXkZZa/huwnr8v
UzhN1O90aYG4qYvmNFBss4LhoNHBklK+s62mYjntO0SktOmW+d61b9Z/4MWUOHAgLaAy3yG4BHbc
ylDrVNXunMQTZph9+iJtr/vUWOc2bfJ19e7+Y1MkSFlRllVaCz3Mkp24InrxsJi9TKpMfKF+CnWd
BQPNyhc3RgU8fOQjMmk0pLgQoefjAZAc9jhjdiMdGf7MInSl8BPkEhhjPuibslm5+2xfYT8qYZ3W
/G5uoDDg3/MBdZ0EKQGqLhxEh7Ee8ro2zQPw2Za/sk862NWClDpIkio3tqL74tDrpiEEcezF4RYq
EJZFYjmRh9P6N+hK2PM7BhZSKA1Slv/GCQ7WXx3+LIHUlay6OYeN0RfcUzdKy8zlD5Hi05Soxtpi
QjtOE79JYWmIZQvQP0Z09M/cnyHrWa4u5WoV2LNNioCTDxq8VXguyKU9nFi5vDLw9DANGkQ+RrpY
ISHaZaMTCu8y5AccwlKC1ma6R+vMqoQZi+OnRlsmXI7HK7Om8E2evq/zkmsEg6nPtrj8xj2U9Gqg
aaFG6rwd4z1QDuAUeRcy5bZEP6AElhnOSa+qwo7kNv3UqGEifIzMrUQHj4ISaVdWrqwe64QxyyMB
CQlt+6zjxtv3qm/Mg8zZsEGfah+H59L7hvecEeJZRVCe6gNdhrnZikuhl8SAUXN3PHZldI8jRm89
3dxLv23IcCi+qloIiOiI2mMClEDWF+efBjjByMYY+xfSGaRZEk7QD9yClNjZQiwHCXDCEaAnCR7Z
PiWlmN+J+jnNIjRqhU8x+wmueBh2X/qLiN4jCf5wACpoZS6aVUNcU++0Ng8i0UlQI25JfA8fZ8jY
hgV2aDdbGMMEK/lMPuX+l7oeyFLk0lyyBuiLPdjEUMohVKD2tCsAWvwqS9SUPI4ragjrtG/+ApBA
tPVaV6STnuuF8+BJ/0b9hz8B2pPFfdENRKkQQiJWVy81S5AZmuTZMrR503WUVFfNVg49GhKOx0G4
61Ly/8oSU4waTbfPhwabVO2UUVD8VRQ+8Rr/J31whANFWpBaZDF4rzbLEHElyP+MdbhAV4bubodF
kKwhfb6ms9wPeYyXWeTcGQiBbmlxxUCjSjUQMk2KOrd9UaND6SNZ1HzbCKvnkihbL4bUnlKlyZKi
UnFhXXaSe3GjnfDAwfaNrmGH7qfIiU06GhznkblWlmjHT4LufAYvW55gXaoHAiN5iazZr/WzMZDz
CNERTz6GSwWcG55jJJOCSKEmYkYfbJYy9l2PIMWm1uMPRbRzKy5j83AjxhbjI9+mX20+VjJ65wwC
YM1+UUVyCur6ZaIFz1wmuFxArPDmopCnBBG7HF3xFGpULaUJbDegzhq2DVwhdV4zmrU/qsPyeBJl
IpL2u9LeHzNcL9RLAlTZpbN5anplkIP9TJ3J9mnaUbQYSiP7oznORRc/dUJ+yXxfddcwhl2GHy1u
x52Q2oUo8cPskbkXL5/vN1/1ypO9aolh+d/e3W1RjMKfrVlAySoAzPfkEKohty2fXWhVkxUTLw2k
XZVEbRdWbuI7FT/8BbIjuKdH3SgK450GI63Z3ANtIIg1h0pnRLcpfzvEqsbsS0FUjawt7FgXuC1l
ZS3C1b31zJuNuZRt7uqld97St2G7/140hPzmrYukPAiTyz0l23TlmWcf8TE07tkzbAKeswY9tF4p
h6Q5KUKMtZhgOhhcqnou2yfI/wR6klpX6OAK5+My/7d89ZiWMpUO3lnCw7l54QwaCELCMdczGkj9
5fAsHZkJTkyALizRMpeK6knvGxBPEbwiHxAz5uVLe06/cad3zJ5esLBmHcMfolILCUC60wMGjM2F
nxhEp/Uyu1/D5KJMbGMaF7L8GUVWddsHtG2g0mIazL3bMbFOBJFUsRkGFF721/o2rn87Z4o6baBY
+Qw8fZckh2rcUOiFWzvS8lIYzlb5xubPSAdGq9VWOaLymrByqe1LEZe2780PaRhwzPzwL23CRYMo
Ok4ig93A2qUhSTN0k0bsLQSyzgSSiHoZB95cqgVu1nFCwuwZuz20EbaL+ho2HenMVi5m5hG4pCAJ
qglz8ap9fiXXwOSwzH7gCJ6RytsrCBTNd+acf2S+mrFfupfbYbshUYrfrEAvBBOpxWQ0DYjADIBt
g7cD/dUDr22V4pOA9Sv6DEBxdlJOUKZr1hj2fBbazwsHwDxs3HuyXCusmXIlVrgdIdKEGWJx2ugH
jYaYvhOevi7XODbKi8vAva5LidVtLNePdTTWrEBOLvfTqStuxzZL3hn9xcoXIAwqQI6N/lYutblA
/FJ6iO6KWyAbonEXB3zn+HRbX1sYeUP9XqkoaD49OJrV4o2j9GyfH/Ty0BC54lrOspbyQ2c88myf
eBWtROE/ILGukeLhmJTSKjo/kqT5SnLvgCG/fEd5Jzd5QGxJhDsSCbygMJYJcr/0GpISCi+zj8TH
meLK7yYXEl828JiobNYycWnOda9WveTZQoIegCVu2b75wItgLfJW259+V+AkktFQApGA9E8NFjdE
xsoDW9Gt/fATu4LZycYIoAtT5f+CB3TBJOJS75OmX2+wBJ48t4/zL8bx8R4TD02PfRB3Wxz+yml5
3nWjl8fHtAffPv0Hdoey/ECPxkKobuNhXs3Q6jiF1aYQItlbPHr+GmZihfSlFM93PBVo8AeRapnP
b6QzpbtVXxBuYUz/4tLTA3v0uFQ4Rxiq3uwbRtaX9eDCxGpBwzJ4X/TEKKWMHgKuC+w0x8+eGDst
Gq49/40nnWUFs/I8+Jm5lKS8s2h0IXx/QYVQnDdA4sDDE0xKu0RSPetTgn7OcbSBYKAIREZdGuxM
aoVLsa2jP96cLJPQjFyuGmt/SdqeU14evFlAEEzgYaJDo8UM87VCP4GkZQX3zOe1V1JeZM666K1x
A/7AQ74y2kBom/lbUReEa8N0Jb0gj1ZHGRemfSKglXDsfTo4UnvYUE5gmwu46caIYf9exxMLhxRP
A/tvLQEVNR/Mabz4UU+B6BeLOwyoNxXFl+vEMfQ9Ic2hOj7tNDfPAv5wD+24Wr7NhvBP61PuthSR
YfHVsQ3lLMaedZ/reS/MZ2XOgryiq/HrsJ8q6x0UmoWKgDh0+WJTVCbvgc4dZAt88z0AI1ruhEVM
79IaFtwHgKgzFJnl77itD5ZgOc1c/CBKu9qb9lGgtxIdnonbmlM48TqvVDYY0Fg/AjQjtH1wsGbQ
TjkDnH52c8ccRdEI30/oIQUoq6cbjvjwYjvXFWPqk3bb7Uj9jUdc7rkK91DHnWFdtiQqVmByds/Y
LmREo9K5kAJDHFg+xCLXRyOJTjMdEcioH+bVEFheH1BK66+gW5tGgU5osVHnWK05Z5vJOyZmBM7R
06sU9O92rGumduMQFpkuJDPWS6B2Mly3P/P55ddLDGlNm2nsFv3HZV2svvFLwahgl6c2yek32R8x
l005Nr9MX3ig6TgAylcpIZxxLGSPHDoRqwEdvbqH36fuIMq92DyD+g5M1vtoTZnI3kgy4MgPTXmA
IPgVGZoMUa42qqrR57ZxXJCKSYL9xINpET3+j9SZV4lKUXBDgIMTOeGoEElzioDOBD2T142Xa6hJ
dPYwV32wGL68I0xOWGeFE/vU6diBH4zxm0AicIRpiar28YcXAIZ/8ikhj640LYTDLF7Jbjkgdhwq
YSWKLlqJwhKe9mljlm6Bm2EUKhmao29sQ0YZcC3kUoBDoWXc1n1sF/sUcGnEqj8Ce+4cLAS3fkx6
GTstkwGzZR2NBPl5HGe8lA52+SaKHLtsXsjF8jMfCCSImxAsjzvcl2B+SM4rYGz5P431UOUfn7LB
WMDno4N7J+ANfmd93QYiX3IQZO/ZqNYOUa3RWv2+CpN8KzvK+p8jKuFYOYk/pehM3b7LVtPvbaeI
nN7ccqPTBihe+mt+robxJvI8WHrP3Bw4iiQ6xxCrH1V8dLW/Q6vAiiETVdIQOdzkgVIvRrSbiuaW
PAsU2H+OtkRDIOB/xr2u9J2SIf7glPTD4zIRK9Cu09t/IgMbaOF3DfYJ+MP21Avv49TW8nM6s2hk
NLs6CxdirIAToPHIp/Gb8NEzs8vOdpYVoX4fM/NineJQzQZ1ZCmbrc610OUTObyzYoHls0NdX1Kr
baYdGv2EQ1hBV+aGB5AB7HNvR+u1zGMiXCfXymyqM2liKruhMdgwU34aYX+8DcxLjjY3pwvE3HPa
R62JE+3NMX24k5by0J+a7VyGsbM482PnxmqdmkhL/9ToRqCzDb3hlC6/9vK2U7ND6K2fu0yVBXJx
4zVWlJV9wp0kNqA9BVEBO+uGncEF87S2+qptlU3X6jE4Peoxe+epdVQC9aKmGd+UXdZffLad7hvt
gdwlRVq51Ti30x3Ff+4iuFidbtpn21h1qXyz3M9MeD0KnMMA+LqAL6saTcGbctIAhAEXFmFYp5K3
4dJprz95lCZjKZRBcTqCUlEQHvYipz4l64sEBNMVmclAeX5/LQVBiDKGl2BjqU7wpwyQWsI8v7l2
yTWNffAU+gFuv01VTe5SCXssT/DlZCAACPDiU32JWaQJMcXk0XuMxvtwUwb8T9071Ku5AduiIJ+B
g9MJLBEgiWAqsJgwyL4JGWXBfA2CaAJpOk+rFF8p/Yk+azkbOV4HmParNgWIeuaDn0217L2KF3tV
GHZQ+oQ6b8LWR+AZ0EzoY21T6g9rj6R4IPCB6RH1ZXIAuOoGmHVhgEveJb2XrVAwzYdMBpzzDdVk
xLocYwcdCqaBXDNjyBh993Yv3/gevO+yW0nunYlW/ZbH+iiRDJPG+Z5/OQ2LVWVS4hgMEd5fSqPL
/VET/6SX70uma9x1qeOQ+ZkBlqoqYvH2pqDtHHy/dkc8IoHD6hogkIsktR0JyfZ+A52ll4oBXS6R
NS86SJWppGPYsv+luNU0Wv5NCupz09GThd5JUMHVSJp44EZqSWUna/1/GH183Nfr4xk+Ecfrlyf4
5ORhp6OEcX+8kxFhXeFmxUwnrIg+GsTArXoY3iXhJnKjEpkElxGFVDl8Uhts+sNyis0qw2smSNwP
pMzouilvtRv4oPpYxhXk6DXFYjZJ3h0Sw5mMaYCpuaiqjz5B3XbQ1bvBPELKcRzg7Cc+d9SZjFQ/
D/Swk30PVVvGFuvOIpdoDVKMerKfAgR3L82wYcZbpYUWun4qqAzAkB/yIsgLo9wzbIeUpJSifnX2
qJ25u0E81XHDFGMxa/rQoIsv6YdOp8Zs2JdlJhIzgSnkjnaGPqgWUOPs5h1eChebuhnQ+zuKfCY/
s5D0prq9x6vv+HBnwAwDSJkgP0l/txrVb45NbUzdLeUPc43XN7a6VfqOpIo3Xe/3sZfrpzbZkq2I
L5nHmWn5nfhXLN37fTUXMmbPqDNnBqx+PJ+7pMfI899J/FRrifOPY57AuT6QxXx9yo8cv+0PYqbU
Oh3+htIgcBwj4e+po3Hne8aa4B5R7ssg9AM5EE/+n0fet4rIiDUCv4RiKya1Korbal2NKLZpdJqC
aLjoDxTVH1rNwIoj2xwwSdXQYJ24bgrSm32ZSup4iKhHOodfRVrwINad0qnZO9UC3DK0Cvntkw0E
12Ir8qH3trrp6+L59x69Oay1kJyUNE91BHZfI7V9sCpKHCsR9l3k4VNOn/rd3oo9NhUodz/qZqHw
6DG3A0kIc+9exARS6J9dJBp6rs4xpT7UBthgDV5XmUmpBAQuG7eYd3hs0Z2o2uDST3XNohNjvLEH
+QtXOesoN6XeCP9z2chBIYjdjVOZ8sjY6W5sQn+DrXGqkTM6jooJ/hvRj8edwxy7xVM8QKbDHwEO
OwezhTsTKTwBxmodTqA39SBAqk2QOUGhUnkbnTcwjmhDWuRx1t4QbgboPlmdHgdtqJWb7thxkoJj
yB80VAD3zHmApUb26b9aZtx5coxtkNVTp7wPpNO8y/Hzz+ZwReeEmkVp8wM092uGi1Gl0Al6KK6K
x/1nVAs1WFfAdgFS7ITI4VTV9l4x54y5O7PiLniMYu8vYxXMVswR1/IWvZREHAH78B1bRPTn6HID
P5KOIRdT6vEqVpJC2bKePxOzGtw3I3oCAeZDvMP6GErb/JSG0WeDzqidj4OSLSaKxII4MAeUW2+Z
06ZNrt9NEBbbrgjmse0OE4+a6lw2cOL1AFgXrlM+0IDcO9WPAp5RtRwue299x8jAWUK+P94k20D4
WLT9jwu9Z52ZEk3PePnfxcaqD3yZd9Oo/An5jyIeqLffqfKNI5HGVaZt1ajdYaZWcX580eHmaPhR
QmDYP5OkaaOSHIbSnqCM7815L8tQcWs9ergs3EuZpF140FqI7tiIvGdclf0Kq4ckbVBq7jMqVwjh
FJLF5KiLJRWWDwDJ9xxJPX0oqIoTgrSk1+hZiQKFPm/UnN/pze2lImyW+zasB6nveGaXqp8M3NLE
nL3vwJuqjCrBkWvCPDvjyfzA0AoA0LygBmQuJYts9Zia50iAH6ad27NrK5AKkUR9CeqElJFUv2dF
fYoG8TG6L3GqRhPt6fF26cYzGwTaYFLRWHSBzp5jZ41mk7Vq1XKLGawbenMYP1s+4d9wVMug1ic9
jZlajlAceByXyNXdbaHpQJMmhEkvPkP7ettWmfKLa6Bh4F+pOLriFs1yAoAxj2uL+g5EvqsN+Le2
ICN9HD9olD9h2KBddlhHR6IFlhAU0Slp9mNqxXtWNJJP/0Mi2pySUMoPf6Kj/lpo0IJsU27+DEDA
53dO+al+VRDfebNEJpCgkQfen3dIISFRsTjmYOxyemBwa9+u4IQRRuZX3xO5+q207WpuHOYn8ZsY
4BW+/uvpsiNgELpaNRWHnM9OjL0WD9qCggZ+u45Tz/5IEHCgIkm3sCmcF2I9w15GzJqyJlLEqzHA
9IEK3KZcx4FFk6OVcy6IUWod34Lo7NFX6R3+KVSUjJ6Y42MAcvKJVH/DvroY5D4S5PNpEMeGeG1T
tXLaZGMMKe5QHbSUjxDTCrD/vm+B2MT7GD6tmvioLiCma63xZlSjT4zkuPxtc5ACAGDR51j2y57C
b65YHuyKCof4hzGWKs8gAQBn3htGYX88aJJehkSupykJAPKMLrwyA8Vq215E8vSJK99jcH99zmq5
9lPG6oVUApn7sKtAmEJfhyLbq06Y6mtstvaEYc1KXBfP28Z7AQRQHOjrJox815jGj1CsJAcpVBWc
tAJefuPqe8DmePot5LvZ+ibRQbb1dPpdw05I9HDQEExUcrPWAcUrVSNkv5MW1yxExg7VyHxrLc2/
ZE32tToM0nFzSdwwbgbSlanb2xVF/h2LRtYzvBRMxpn/j4zotb6E8WEfN+C7VUJwaZitONbiPJEK
Pzw++k3gWF8lrQaoA3N9SPzzHXZWBloVTpGMCPlD0I4jZGK6TmoBK0GOzaR+8eKyh1gs110hkLF0
hAharN2EcuR64iKvYtwOgZ+PcDYDIzSmcaFRVO7ke9GWNw2IpbFhbmkn/mG8sVTSmOR49ssKpNqL
8XMuHoN5xXVoQarzY6Rj9pfAGBJWykYk2k85tuC/WQgKkOhKJDjEKDLv5Ikm8vZ6X+ds+MvEsmk4
jttKhnR2N/l0SvkANqqt1FJdkWJt1d5qBBdgCFKwY4YKuIrfquyMqiKbHEtBbon8Em57RDrA0YsX
+t6LS+XjnikR/FCjrTd/pJYYx/xSeczz4nmrd9RdhRsEKFoZsClMDU10z1OaNx8znuZ7LW0KOMQb
1AqG7mWoKIQrMzeYxqv7hdaovxMP9GDj5rbK2krY9TBbf0VJLqzd211++ZvUKwcYBuxDnFN7c43v
oOh+cUDv6ehnlijXRS1xKSZ2zR1xRfNnwHDjJ12n31rLHzWLBHs0TZ2ZM4sJOaRIk96Xk0cYhdTI
eIktkRNQBv0KhLOMRVUl/mKf9THHRKOuQ2cfbt0OgbgoIXaaJJKRj9gEbqjxk2oE8u3qLuLfOwKf
IW/0sjgsyz4DBWofMirvSI4oYPooP0FLb7LlXu9qXBoD0Fc7VgDU0vMVvPwj0CxN7IZjMQHgJqtQ
tKBbDeZYxebnmROJQboVo85NCdWg6UKonZmuOf3/AeASrjiwTfyz3TJ/dEaoxB9Kf2/80VYtRnXB
C8vqiuaaAKBcHEGkQYXYoViiIbkgalgVTHh4acw29klEN32a2iS3cHgyjhWhQAD/B1Y2JuVfaDCg
hPEzf3KkAbG9buUTtPITkCK3SN9W+CvJFiiafPa1z6h6VOq+ji1B5PWSA3izqId39MR8h7mJQudf
gQY6+hcWCIsSebDRuhm3m8rrmztaqDI4YIk/CLPBzQhslPEWm0Dpya+FPBT7OfvuxJ7QsROK+XSX
1sXiFRoRPbWr73CDvIrhfx/48eIX0CorD2pURFmgCP3Py1avM/3RdCF8PjeJSsZufHLs1VWbxH+l
GjRNokdwgPkiDDs66BhSnmhk1GddUwfvQIOegiTQuEnSu0XGHW/KlnhmrdYR6GGXJa95Ug0C/qZo
ihEXanvz3KtFumNUSYhFJGe2+x97q+mDX5Os/LnknIYL1wcin5iPidO0KaxcIURicvA8o6bQoIRi
NQDNnjGImciPvQ7Ynm3FloYzVwcvls520Oq6X3lGWM554UIAVLZI87UGXR4dOYX4FvI2Bu/fKlZp
s3c7WEmJ5gQbcKN4f9FhPHKBRuuX+JA4fZ4FZDPwYnn1FqWXwNMBkch7NttTiLFJVPf/+LdMU/iI
KVnZ67Uy8bxHepTqgTZID1sXDaUmII19nthfyF5UQb3ESzYR7D6Ylbni8sjlec2ulwJwJCIOd1IL
0JqCiAt7FikaUVuzqlxpbP4yboIW6aYtrmbtibU/Zarna0CF2jGXqMBuEu2CtibHv1zSMZlCutbl
kSssPJAnknxs+NGK9xKpA1WNAlVmJBD3aH2GMRL8QUXTs+gsgYg7nSOzaTIo4rstG6mC5jgAFlVy
+eOHcRNRIZURnvO6k9gzOD0CvkP7i+SuOwIEc/eByqOetWE2x5Q5/qvnRB7jbkjYEUDUzgvpsej7
d/HtukYzPBOr1yDQsiXFwD0//xBRqy5slOpXPzuktr/PjUGYlNcWMl2gmjnhjC1Lhtf0K7Vix7nF
Sq1Y89e9HmI02DIghv4vFfO7ZQzwPV3u8nNuBADRLt4tqsN6uPoRm+NiKuYMBly4QKxlamZLqcAr
1VnP+/E4NffMUHBZOC+BaNhiOw1Szk4EEkPCu6P+WbXkfYIKodmTIBhrhy5mCG8BVvNkyUTI1B8B
8lxNPmTUQPUXqm/BKvp9a0PdVt40CW3y9hx4NDg0RBawx4srtcyOsUoUMCtUSwa2a9ZuEOq+P/lK
SPs1ClPdo3Jg09KlDZjU5vvJ3Xudg8lFZ4pd+unZHnLxRS9JafG+9vfjQl3U1FOThS8cJMn2HkqM
p026a8QmazEUq1VZfCQqjeGVhnLWzNYzpC7HyrS57bJHTeOiRws6TN0Bktn6uVI7pHKilmqDSCd1
lZJTMuFdZkyIwt6bluGFEYF0gOD8KctPvfCkvn8rJwuJvqJixUnvpYFqm5115sOH7jDZiNR2nZQe
qINfldUy/jkwZUY94eTOQxuEtpDLJDU2nXqVQhAog1dXjoMfLzXuFB4a27RDp5zuAbDznDtwXN2u
lk8e+mvWd46mNLyDbnXpFQesbTwLSwZo7Vi+PNud+VG3pYEt4MXy5ZEpMMHkPjWGBWNOc+XAakpC
5j5w6C4spUy4feP2RCGCk8zlEi+1g+kgOxx7Y6mdr7PBl+ZxllP8SY5pIYJkc23Edhoo+09BlLpW
bwCRL2VN7TrkEcgl6VhtjpPFGddbgmLxi8uQU1GuhmwMgDzb6oe5VJ4BkkwDZJMq4HEM2EzlZ7Bp
Q6mN84uzB95IWRRRVOQVyrVfLyeUOTLfNh5KM5FUaQ6IoYbf3k3yhKGjSajPogiFzeh2ggiWSvJr
krfCjhjynM6mmk1iztXcX92jx+NuoVMBDUoQVFN3LFGlBEdAhqD5iw5mEkB3C7JQ4OTYkWCVpmOk
ilV4evejgCl43O0BWjeKn1vp1tCcIJL81ESg6/BV/yZ7pnCOg8tVWyRQgZoX3xqvdJqCAM0pjRTU
owumlq0kDeI1sFO8f77oH9E53Sy6UKTfevria+fS6O2z3KA/rMbOz9Ytrlew7EKFUwN6FoZOhJB5
qYTFJ9g6Y91xn+WnQ2Uf1QvTFP6QQsF3pLXXjd455crNwAy7oMj1klhMVtY6S5lmOKrxHHfAi7jN
Kg9Wv+FGNyBOCdQ+Vo+GtV2t76I3roLOGLp4QxXLG9bPpPQ3hx3BM1+0rJaM6BJba0bXksxM/7wd
ipquwfUPZa5Yg4jC4h5jgZhRIZ6Gcf0Y7Xxk6hkdT+UVrS7TnTwoFcd3gyWJ91Q88FN3S8hENC7Z
VTWNIUvLA7JDIkrsfIgZonWzN3rZ/auzD7aco+tiUkubmqwgnfXfUqvqbcp1yaG7pkiO9jy3jrEI
DrFZTTBbiHX2G0KK5Zb/h8OaFfBln4hgDpY8Zlc47TDb2hMAsLUT/uSopfaErC3mZr2BNGt1kSRM
F0Dg+6jw5Gvlf4RKjJraF4hzOpP5n2pyrp8PD2ZkAyzpJogf6sE3QmZuDXOwgFE+Kv5+py/xQXgu
ewJH1Yo3sjlYLxBE2xNOtTpKDQ00rned6aiS5ihlxXUp72qyBMi2RYJWLzcuIc726Hhyl92FpbqF
8nXFzvkI2dxO3GEnETrsgaW/Eijlq/t+p3yq5rYJZ0IRerd3OVHJnRVmxfwkiL5dqtYcaqPUcmdg
Wu2DGnqPNJvPiuo1n41kbPYoCUB+L5yN0JrKtpoHTxocNsfNOvSYHynSADuEnBaJeHzrIGUlQ14j
uumk5Scrx9v+KLvkWgBppbsE6KKVP104/8FmlP6Jys3oQeZJ1oTIUJZTEmtsnstXVHfAf3Ab6e+X
ZgKMA+f25ue8cL4byvPFhxl2+RBTpc2ebpO3Kj/ixy0fOQALlLJiv33NIvECug/BnCcUw//P2fFl
p1WrnV5Q03ITS+fU47FswJMguGYSEcf6/+/F3Y6pSdmzzz88CYMVcmPY8BtzXQ0OxvvPNACD3mUe
YUBHIqJDn8FM9wbfg2ZiTVR7N26cLkwYNZ+C1m3o9hpC1Q128QrKyHVOCb60wecbsPlxQ35raFMo
ZQk9ce8nzIFs4nDS1551uNBcL4LABqVD+IQ3nPYvQaMzV+JGm/GHZ29qLSTjieFMujYxlL+sqr2Q
5QkDXdUQ+We+QR8y5hdUJGLYZxv9HcIa31fSBR1va0zr7R+kE8miPwNfiTtfyUOo+KS044I4u3mg
tOPe0rN2LkY5NZL/PsVsY6gEVMob6W+/tHhwBjELYyMSoELPKuuM35/YY02gkVGe2krYe9xljfsb
w7ZUZDNQkeUN3DZVZrkr7WVmoeUUox385fX7wcrrOoBk36n3p4fx/AYlgK0o0HlYzqOuA1DRLMOt
b2gJdYaUb+n/ObTBP4EUvjlXIQRws39+LsSzLvUzNhyR/EAQbAZLL0K2JiPU9mgsJxqzUuBRyPdN
WYfLUf+GkhPK5AqR6kjEK8ybnMf5pXIopjEeDCgE1vtHbGNRYt6MnM5zhOEfUf18hjP6/J0T9HMU
2n7ycrAcSAhTvw0HmTZFgC7aPZjoehd4zPYTENOLUDaHn3Ie4LPoL6HHlxjfgOO05JdJEAI0KAai
nfcpfNii4deVN2yJM9ErB2nJcBWOCEpiJZ36eMYtcgSqIlMlgrSm3b6//jA5ap3tU+TM74EyNC1+
2V67Z+WQJ86gbSKpyzDNSU34SksqKbse5zBOtzWmWMovsPNrNsQEkfna8JPx9AfJxCE5MUGN70Lc
xj3Zc+i1Tdur5LZKJEf/aPUX9agNJogp/eYJoHbZaG8QNij3bUv8+yoaMFHK+GJnVX53/SsZostn
5l1hFLpUnqg/OpNJ6jdPsm1nbrB9AOKA78UKMPf3P9xnJ+CEnb5pgzJoOfsuvA6NdhAGT5/1pQmO
t7Th/gIHX30+VLFmlK+H1zRbr1fZHB68W5oTA08qrW9ak1Bb1hzIdhtaO6Dtm8UARQb46+/lKRHY
fDvEsZWpvidLqs/A2iKenT/R1ZyPfAVm3MUWquWf2Zf4Gb3DNQGuMV+yKv95OHqF7oVw9xxEuX6F
T4ZPyi91N8l8aJPz2ghwyaMmw7ij9xvQdjlu0agxg0Uaf2N0xQphxziTannMiBblH864sJf3kXml
hMIWpmDscnkdz2qcPw0R5LkI5QkaSUsnaS1eZcpsLhRwO58d3n6efUW8FxUZNbwIzH8achPnKEAC
ykiyj6qliVKasMAtDDzVhif+kwECadM3xEpp4mYowuHxAs+zOfQh330U591Vn8BLOP3M8OC7U9/R
JS3SdP7c0KEBfFCvShqTUSBxH/rtBM44YxVQMYfh5fJESi764+9SmPQDDr+mT78jMNJI5YRPj70b
Z5QOew+9SO56HWFf0Kugj9TdB+8mHKIPZvwG6xZSKNtKVe6H2dPqlf+KbarG9P41SjwIYn68Pm48
Q/SyLpXgpySTeH4bCSj/Q0SUHLXiSntWjWPjcP6iZqRjD/yibZjIvvR7zZ8k4JvFJ73NgCinNjyG
2df2Y2G9VQ3DvFkQPo3iAUpIz88oWD1BV/SNJq4tfEP7P1fqgWVg09zA/6kYNH2lzfPbw2Iwi71Y
NI+D29Mu5j1oUizQxIyjBICXwwzfIo3qpezi4VCoY1y7tQZcpM9+UeGJmCWXrp7yi0i1s23nDewf
LzL0Z4C+JTziVv7Wxw7bTPw6ZfPQYO8bebMaVo+AH2kZGRxA+sRrPZc+UOv2z4vjAEedTw1yCL95
hlpRJhuYe9k39Kb8UY0hgwGBAuSiuhapMVOAlNaDNNhkK3ODjDvkjWenjg2kqas4d0yWt7uNoIYD
FBTcFuiIsdF1L3kK2i4It/us7OGeZ2fLaV/WJ1WvEh/V0gxVpjlkdaD3TQ40/kpGzdPr4CYA8OWO
wl9qSkxa4G2L+8e7cUIEmvgx0nciQzC7f38zA92Zp81MWyfYecUpYh4DoxZ6MjB+hCrGthObEJd9
LPs9yVKHr7wZ3U5tg2wp13wwqfJ9YjP6a4FC4YhwWJVybv+UPA7n2xe6XFeaR0B7nKwcFuhTVCUf
OxMEuY+tJvL6GeU6aRNaioOCNprLTXretGkXLV+I7Ssg/OgsY/zBAfJSf5531SkwQIyHDHYHu3xI
Co3ZGGg1kB5wIxwJDCupBesdkv6z7eSfsytlcgxVsNYdqWdFnviuFBEiU464j42GMVpk3yXFB2YV
0AmYPT5G/jCCGIILvxPKFPdunR47BanG3fBbuxTX1RVv4ziHiz1zuMvUJu7buHxYH84zgAlC/4PI
F/V781A02umsT8HmcmVnI32CzxthwIMjChxGjaJLMou+yycLXhB2H/kOGMihOxzXX5oowQPRnzla
ih3VV4VLRIfsb2jU9YO6CS7NtcorkBdhGKo3nHEjsyDqdAheYUHdw1BMb5kzmEBJxQBvQRN2m5me
/kPHyuNerAnItnQ8IJGKFKeUK+MNy4J88UD4+Dlhd8aCTL1I1zFdOhytHv4OCOuDKVWncwP1keBa
TnswEjxUV3uqndbxIcw996xt681VdSc+KneQUW//rThPfowZRow35jA1zQzkJy55kbzZM0j4o3O5
sYvo3hxGFHrCwKnnymsDM5xBcPdtkHAtRPUh60YRCdutQ7qbLxfptESBRgUICKzx8EIAtbZZIEKt
Dx23W/lmiU5a7OPl9f8a0D16ZlqrPJ/l8prEV7oP0lo6MZkb5IVkpaqA4kdgkEZVs2G+zcp65uhU
NpbG9VxCEXG6Wq4gB5ovqtWreWjgqerrKGYW51dbHiiClRRqj7+mUYxJsAUi7Ub3MgbrE/LjFJBW
Zf7wouCc1NHezKEP+deqI31zCML3xBAKjbJPYKSMHQrA8kdaWJHp17k/bjAdmAhIo/3JLWs48pUC
CRenwsRcGB79+8LT1jNmR23scl7zjcX8A8WeILGkd7Ahk07PeMIAjXfWZJsEnsLY27g9mD9c6ZTs
cKJBs73ahkpNT/SNi1ITyo5tCDMV9HZlCuOjvnUqjVABl8jMWU2S3RQxUc6FDG5Nj7YCIVR7zYEk
4PsriXwkrj3fIrNYBHRei+ON/vF3+I8cN4QBW18Xlr0ImV7esmR6ouQnbNGgI1vQI3HHzGsXHbi6
tsSSAspdTwFWaRRGFxE0PBVwpzIxSRWNxZmaGQgWaf0jJzLsCLK8hK403T/906Lrbj7vlk+38dXO
80GHO38lAFf0LKjlAZvIsABeeWOhq1KCSAH38rf5BfKaOO68R8NJDY5fA6IYrTCv8bPI+lcXYC8E
n8s8VpzICUKmHHypT8umFTesq9uBdp1y4kvwyXHP5fjMnSl9ivcG9MDC+4k6MkQqg/Mfpmv9nmUn
qykro3+9G/YWQDBISXT5xuOMCT0tYqSIDEwzJ1oKgox7yqkl3eVKvFMsAn5PWPGLwyUXQJFUTQ+j
lcQ/61YJm5pqwRtbbdJOmxaOIgkdtQTvuZuwFCVc/yR5iPWH25I6oQEIzPJmbcBCXsQtZ8s+06ni
tc2orvI2fyQ/8JrWXrquGOD2w0fmJjWFpdVKihsyyR7Tfv46woaPk0G8YfCgUNIB4nZ/xcui66W6
W9JkeCJTCKhkSWeAD/VXHpUylUw2qJYzNtNZYKiD5sWGKlJwwnWBiAsfeviwjzbPh0g4nh5VOyWb
XzOE3lyXlGgYB+3oWE0mB6p7TjQLSwdUb9x4LAps3SGHtJLIHNjmQP1g5Pp6BbW6cp/fcwx8gpjV
r5xULarjKZs0OMYtJ5gAY3fN9tXULdoZcnVJMzzB7WW7YLsy/EbNt2P02aNaYzv75QkeD3Ctlejj
rhkP/UlDkAwXuYb6KSVaruOTjivF0RVOPcxa5AHIWnUs6r9a9idG4HUYIprZVvMZBqUcf0NYPeIA
BVglNcXVUx1Gk3lb2/lFHbYJ4HsgbDgOUGeV5SwrtDlChp4DUqFEh+zowgAyIInIkxMcFSp0IqMe
HC2RYX7ePq/QRaYpfUj2aNd9QTO+3zRFWO9Ktt38n51GCU+HA+zxVyQLoH3F11ryv5AsoNs78HYy
aVOMfzSunI8u8qOkDoD20j4UdmrEHVk7kD/2LV1GGMg8/942eKbxewXF4ODZJOZr9ZQjP0lHTLml
9Ce9Jh/q4ygU1HcYVCNvoek/uOfh88EBVD8pmmrYMnOCqJU+e3ZbKcshak7h9rUqYW35hvEKSpSs
9eFZTXve9UK3adJAt2AjRjD2+RSPiEoGvq9cYJmcrnifpz05ub+4IWaW+JfCfFJfCshIlTOUtgIu
M/lggOaIs1AcH+nvg5lC8tiQH+3vZY2tZH59CKbViQDgRSjemdLqJI1SxMuWr5cWBs3rVrL8z235
+2OAgGoG9Xk5SOqhdrAtKfqKLDCSVaICgGLx2uVykfox+bhe0R6nLxmqchYDalCpIpix9kgMXWwZ
4HrV3vfFvxPWQwD3g1YCgZKRnxWDMtwkag24pnoRdRKnACUXiY0eeNFGeGOnA078bVhfgl7dd4sV
cUd6qdOycRe1X1auyrX2VhYf4X5UO1cp0ecCG5+WAUfgvFiMGggT8Rh1107+/QkHfdnt0waYQl2k
t6XARCz0A4t2CQOk+zPFpmWUtlES1xYITy0QaYT7GEY7tPdIRfKS6oIjVU1euiKSFSuCirNiAxfZ
AmsVlR10ydsYS9tSTiQsmoURFPdin1i+lw/SfDbwUf1L+YqVHlmw48HuhkJZ4LxS9Ekfzkov5ng4
queREC/G2tAwaNPSO+1Nw5GFr4Dn80xAPryTe5ucGM4qYSclKU2tGuxyxtLKpOgi/1R2+zFJi0vD
RrsCNB5H7V4PYRcHw0YmlMGtztwHSPmwfDtbcLNm3uS9GY+uE3x5qRMsjclRdbxqIOeX1nbzeLsF
wW9Shht/XcNJ/2GAkKv1BqvA7x6dEO7k3ZYDGga+1/25ugASvf+Mpcy50ySW2krffLnaJ+ugSNwr
9hEs/cA5CT5lbYeP142Ugw8dkIvKoCDe5dXqUETQMVhk+sisSBMLcreGKDQ6fPwChz3tsw8sybUz
G8/LWHhYjyWsDmvWmQQ2mH6w1fyMBkpfMiZgZ+h9jPzAV7K2maz2fGiD3qlDJoMyg3ceCenUbSk8
MNHg+q7wEpKJXlxgGqzJYorsB2hZB2a6p1NgOjrYl+XhQPXfcvrERCQGRbpmc2g4/5hMRd9qLnZL
EzorY1CCt+x2hjePQTECT0Vt7UjMrMJPvv6cizCLzAOV3b8vnQrC7K8dVdoHoGw9GkofU45fvVJv
H+d+V9rXfq4AX1NzWunIRcUDVhmd9nRRpsJVS1z2aFfoHaiHjjY7MEXCYSM9aNb1YxaGL0PspLtR
ib5MkCaNJ2jQ3VYrGLnhhrWPfxASI9dhKGk426f7plKst1puZZAFHLva5yCvr+vTvXntRN9Y1AGL
Amc5Lh9n7nWpK6BkwHMl1/KY+T2A2TONI+5dpWDTlEhymjPnwfSNDI+2LpfHml+FBC2X6A/DU3kz
bxWIkwr+TMb+DOko99EhhVVeIeABOuh03ruyKQXumIYUUevjpO77O0pCkYgTDDEyun54Hdni9ylv
01y1cTWc4WFYIrjt42YXQ9u9MVWtOVybzuIuZjCKJrcbGbeSl3VeYlgF5X7cijj1rcfNKrbUvAvf
5+Mf+c8vIyzukkA/6B5+H1boahHHqdpeBTbcuqBKZoV540QGGRJ0f0myKKwMp+Xg+9jOjRteM+Tz
4KwrS8abB+SPOrCZSXT4fGPj8eIcvF68KJuBXwd15IzOmsnpPaJqbHR4rL97JYJGxn0Aef2mf0ud
9Sjud9YSZ5676UGlr0FZm21/PNME01U2NAwe+e4YaseAj+w6XhQwHxAXiKyNoiOrD+B+ZNfbIGhF
e45eI2GuOeNWaihG9NjOpTvRIWn+I1bib3mqr3eaHzMAL4tbojzQLOlK0Q23pwbdMFzphFRmJxTe
DdIciicQDS6wOjXKMY80vGlwXcBxeSVpLnTiEk+h4Pkocnp04wGFsyFY/zJkTbihrI1BZPNY46vg
Jy1gZRbbVoMEVDxIxn9KpPmZojjuUQQ7djSzuVwEF0pyMrGvPKNVY3NuRWfEQu5HQBHcbzlWCcci
ElS6/j8QEF/AFdlIX6eTrYRMY2CI07+8nREcmTEq0dei9Tnz/ixtmG6FN8y52r7K/yZ99cQczM8r
FzT7hNGR/+DecNxMsXyJOYKepzJQ6OEpgxGilPO8muY4D9snsnHQM80TrTMAHe2Gy6WBow1ueIER
TTjwQ838HguxpaJn5bcBFQ3PY0SFF5PWNPZOtjFyYYV34pl4zZkxw0SqLWoEYIbQNSk0h/rLy9ta
0ygwEqVWn1lXt8WADBalzkOt1lOOIz+AO8SKvc558RCyk16LP5kF4cUz7hHb9loqoGC/Q7eetNi9
JNfnRFMhvME3J6rvsBPPKpkmyNxYQf0rFn5+nRum7sgwRI/oiz03xWQH2OUA1E6EJKGMYTnPh1gr
ePFBA3bOJXnWNurI9j1za7R5JFSTV60QW7FbSb0YLTDJOfpD+uwj3YuYN4QqrFhKSX/Vcq6CDDLN
m3WVk1Lwxri/wCRBshWRR3O4WI7L3Z1kCFvMu1im5kdr9oXq97PLbtVyB97cNGwt3hDEyt3OxPms
ejBDsrZ/xKhL762JeCQ/HaFQyWp7ZlQZfvAwaynuwsXyBCTgIzIEMagihg1Q+FLcjd5kmHOWZicM
KWglzxOAdRt1/MFT4BM/Q6UwIged3DflT2xQTUTqBXjAexsItaDWBpWjHj+8zwdxUaxk2hEWlbV+
sB+76iyY7tA/i4j3qQkmEuS+yeuRS0J1DFnuccYez3oIU89fXZeYv8AR5ocgPPezU7OmaBzqdDOe
LjXC1Wue+H2UMmzGI9YRVhDTsIDVwlzaHubmn9VE1cJBBZp6l5jKfP4waI/P6iuHY9M3wAiuTtZv
7fTzvDKAnmjPI27WHuZLjHRuf0MJ7QCkfMbZVqpQ2wKmCYUTDei5KkHlt1FYaGcY+GtK9GSYirKO
5WKBQJO4fbGDOmbd8ehhjbI2oEZof2TjK9z9F2ctcYyFFXm4LgkdVcqItvfrRTxQvq8wqGkv/8+U
8NoDf8SVBsMM6HGVdK1keG6gNj7iY5sv+NXrZbX6iKYPh6x9PzpGV/jTwjrZ9R69IhCzXWGw477q
P3gROYlBUC4ZeyKO0ztaFp0qiUZTeycDCOLYkqGdxitWLXQCWoVipeFZLYm34Ele4Kziq0QRc9KK
0pOfEv2+QdOcE0xpdI/R6fyBAnNQwtwWbYRt0X6nV0VNvbJjr0lMZWDRagJIqIZJSDS0naUujx/b
2qfFdKeUW0ynAOpEqyyu4b5bT1KjKUa2KzHTKh4CJfFELZYIHuBqWy+PbxAdVGKFVMqvGu7JnmRE
tlGN9NVffsc1dbff3CBHGGCR8AecNDO4mzR1pTgWJu+D3COi1Itg/ISIF5+nWZi45i14XxQL0dhr
Rsek9wkckDOyQROGZ8LwiphEUSPGQHESPSvZRgCFAonP1SpUGmR68hc8pEB2FjfWcqiCp41Vaaju
U/qiJaD/paBtN828hg9JsFtUg7H+zCggTC9qpMNm9MkaJsR2O/I518OVs30wcy7DgNBgO7zlvyXP
v2I9gpCwI3XJ0jDOg9TmnLin8p/ld491Vu7Bph5kldDLIQPTDINxDY5UZO6bo4c3pBuG7Q7ZLAOD
vvqV7J90q415GObU8CPAtkN9HIrhTQLEBL8vl2Ih5PA3yYHQMrFoZv4BNgUKefYTmYQv4oTMQKnW
aXCmn8KXp+yLEfo3NlxFSOzGuEv1kioK+WROuH/IcEE6PENEJ2ZPRTbNDEzWzUNvg4N8J/1w7fof
0LSKGPX7SxLUEwC1uS8SzSsfPk7Uh0YtMY6nXmFYbwRAM5wTiquswNGkRsH80eZs4yPGczRixx+C
VlDjx/I/kg5NDGvl4V34PPYMRr8UXASBFb6aWMQ5zu8zF7rcgRnyU+HmYgqN5HKqdOW/PxdClGQ7
ymWl/sGPddmAtn/tD2/QLvrXi3QMOnej0C9q49KZ5c1JFsfpqctNHKQs1MIlCY4Gzi1BUjzLGYaT
ODHBkeVDxNOGCKQ4M72397r/fgpoaL3CkhuA+P7fM037w1feOXk6qJhogpFOj80FpGAhdlV470K/
DLP7nquqaKNRX50LZJoqHVeWBDLTJzB+FfbAOy8Tp+yyvDvMAdl2+5CUjyiKnEulT2wIgquSacoR
jVs3vkPCXIXwMvCed4V7FdRQnzPkQdtSohs03JQ/Qqe/1xQX3dcU2OFuHguryPIhot0jTjkKaMN8
NddpmveXjzMaIwHkXxb1/Z33NF5Ns8M7e5CIj3NThqPmi5nNSvu6cA1XjkS8x5Z8xnbDRvsWluCF
BL06KOQc5r60oi6L9KoFEQdOXXwmxidn41uijUq47pjOQuztnuASLPrYyXI8jSg3ftRl8hEKXaG/
JBj85m8VM8jkNym4t3AegvdfR8BHM5kXi43oqE8nUBYtS/mRVVc4xI/SMf5PAmfd6Xbg5B7idBlv
Fv1Uf10b6/1o/sefXHNxmBNnUHhypYqma/pj+inqUSSI6XPenGh7aDyYKFr6qD1L5XsZHrKzZ2xR
8r/RHNCT9v8+75FrQSYrWGcKbwGlPF18EYEtwQssEZ9SMwOXgDWZvQ11y3Jpb08vAQWVypEKtu5e
wTAvvtI5rOIomaQL8cgbN0c5fTO8r9HgSUCxFIjDQ5FLxVWZp3H83VtJqA4RUmkh8RMnR1flPc0E
Vwde7bhzZSt9A0Cwmw0UIjSv8LSVmJX37mMhv2Cj2fUk4hsOeK9oMiCsdWOdtBZS1lD+NvVTq/KC
5ZdW7qKs0/tZKewjCeFRKHApMpPd+uUtGNJQALPQA7LiH/h4ndNt/oDN/A4TnbHeR3MixAD4Ddgv
0kwqRoku2351+ringH6UQjfE7qEw52uzk1P8xOJh5dmWvUZWHrr5KMmkcF+OWvQbRyAXKPCvk61K
mS+yaKt1yiwbUKNAO9gwW03lusKDPcyQMPBVKMndlKPfnF9ff3h4QkL4ek6cPUprbV8G/G7jZWb/
sOiFZItQ0S2xBZd48Mf2puzsMixaw5q+TWLPaO55dw0BmCMgt0OHsPuhbxFJ8asnXATYNOYeOaOr
c9nvCJbMHJq8BCQ4AaO3cZOVZn6GfEV0TM3KMCXkDiy5R8aH77Zf6Es3696lxWsuU3J1tbtisYPK
w5kcbShszgYsdIpAWQmYituEvbcngY2DuKi8tC/O1MXRpfvZsE+5r896nKgbM1k33Msft/ZY0oQS
BijPzYYt4drqzA9QpD/G/mD08EMmaJWBuc1el5AoAMI+0MrRcHbQGtpwk11q/qlUcISKQXVOmGeR
kkvMLVNkDTI+bPYftd16A8MsmYFataN4rm2J4HNivRIZZH00mgY4toJrG6WeJGX4eJMQmMBYi9Cp
Potnk+gWtMrk1U9MlI2ISILSj9/1pSadhAAdlshM7SPW6sV5uTyEz9Y4lUSETwpjeWYpzQDcCUC0
UtOxakc6+nG8oVlGBdC74Z4KoT1BmlSfE/KQnQK4oS8ObitcRRaoy5J96B2cO7+PRCyqNMlZQQeQ
wAxBcefFWOBOl+TlvaWmHgDXDLHUv42JRHqJ22nAZ/R7wogQ4NqVSiUr4nA/7voxgBxoR0hD3ZAa
7REXyMIUzcHIkT6PKUPKl12Lt1Elv8EmCBcTie+PZ8LjzT5qagR/V4T/M/UJNAbVkzoTOmkhjThh
ir3h/OLY26pTZZ18iMNzVkLgJ0z/TvwqAOfsBjvbxxukJXABpLSiRRyvXWAS5bdacSwzpnDLOutb
CrkdgkANjpDm5vwlMu2TExDNOMbRYAPCnHrT4Gd8nBRCM0LwpXsMaoomkimBXtC7XYvVPb4iFZng
BFUnkMk0rVCCZ+Rejt234j4UYlmnGZybmT5iF8h4V67iDzPqY9rSLHIIQRf6rCO0KM+Qw+4KgZAT
xjCXN/sVPQgTaDgSKVBoiB53nHoATUlJJK1OEGF2XhffOQV9tHme0FTi2UdAeNZ/XY5XMAP8G3tD
fmqMFLrUv7q4T8lcrrDwcwAA5tCp2nOSsQ0zTc+mk20ryLJ0brffZQC0DOrvY4OrykN0QeIJFqqO
aFuDb7h4948Mwi8/4CBzp6o2wWQIFt8kPN9dpKZ+E7O7DnbZOdHi+0pBUof3tqNAvDhu0DlH1kWg
ATLSZovHGPvyx/ndeKoz9L+K0IAW6/BQaY5b3C+otCmt/dG52V/tZoNmlcgmxNhoVBkFSe4ZOIkZ
OaMaZIEZrfMVHFZK/FZKQwTIzB7uKBn4vyJ+TJQOx2IkZzH2+DCj5ShfCgQQT6hFKZSR5s5znQdV
3YFEe3ZAPKXKB+FJmsLsrgDFc4REQ2NJ2CfGX+TMSKxbBn/caClELmREl7t59PB8NPxO8jUTh3u3
rWHbHXrrOgKBj+GeEq0GYeiO1afD+OLn8LSpJyM3C1Upj3AHLAwWe2mm6+hJkn6jIOI4S8jZOvci
O2mNlCywbRsF6dj0yvwwJ5203Ecjv4QgJ34a1TJbIj6PCyGTXAx5RN3y939tNblMNtDJgagZv3Ft
zyn9EDSYhmH50C0uquR4thnmwJTukDB8oxQjsHihe/SHnmlJ/MGRDNbqdxr0qN1Hbq9w9/j+rahZ
4XZfXGJqUUZvhNbVm6jmo2eZgL8s5aNfx0MTIV2FNjz/OQvD+Zz0fdZKTQvHvtKf4NL5QSZY8+wH
AyqvoFIb4putdXAH3hJ18K8q9umM7naspZ4qdv5ENz4LAY+6NXgTz3uGvhMLzt6640+Do72qsaun
pzhSzC+wM5jmnpBgsY6ehvhsHCOO1WPYNUm4Upl2ek5EN5Bub6Wrhi/wElHtuw22UJ29jtnORSos
+QU0oHEEmpV7kLB73+wMxVeh9rWXypSOKBUdRj/HaDel2gBSGsqkdEAXp2ImuN7cIgW0a4patSUD
UeE3oCGTG7eAGSQsuLQYE1Tmkv8NFsvefnx8fnht3HdRfGSU67/tL6KchTkBna8x9FJ9iyF8rp9P
jdAnHU7cQSGQese+GA6VKgM89YWtK1mRKPpN0kfLeIrq8zXCnDez4nHSZfmD7bBiaRhgSs3eljiA
mBtz+J0rd1Jrf89TX73oFU6gMDvi20ppU+Ym/JPF51nksdJ9uAGfkHvZuzlfFMlE4ifHGNqeLEpA
oo+g+/vdISDh2/FmTAqokOWemxTiQDX3GjQ3icdVOXoIFlgMMlGyq9jtrx7GL00XV3fRaMg3QLy7
szcwuXRYuuuvpCcvtiqmV0Eqd0QC4u1kq0kdRysqYtEBt1pT75W5uAsJeyajcVxN9papqpNOWTnM
u2a6/TM2nVhcfIDQ8nTiJoSr2u+TISlokoVjsssCazQEjqP2V0ghWcQGeNRpybmcqlfe8XAMZUNI
0Cd1YM5gPjaQsvpJHUOCBc+rvCkTzOv90PmJys+I6jwWb4E+GcCMm95XCuxC6grxyulFXrXlPweF
l51EEzdQjp5d+g5WVveKYmouorkCs4XVVq4hVmEuRwLxwdgNsjV0DXbhcrlIZbhj7Y+zKYiepXOx
xwxYDDP6fOryKcSWv5Nyrrs1rdwIG9bDEJZ9enlByZMoFYqfuiNqbK/nDToO36vXJl1vFZyXOrJt
jlTcsLbqajCLWRL5Y8nf0AlXM4yWG73R9/ka459FrfgYQIDuheLr9WJ3ltrVepH9M/NwTPi7lDJp
BKMGYhjSM2ld9ATRY38GUUvig5mkSnXaef2gwLpf4T99lMpaFPxxy8ihOuH4P9ydcL/NCt27d3/u
277yDnRxWoTfCSJjor8H4NfAVsk6ry/SzBEUvtrP4VjQoHVNPm0uGa4kNxpqWLs5mQQvOfV/ZF9k
BWngbonYowSVTGbNKHP7Uu8nzr+/QQvzZdrv9XsOYg4xrMu+P/0u1/rTFUX6SuTcPKoGNweLg9jz
Tl7X5Z5FVWdBp7wb5tx0v9xdoySqHGcFrlQMCH7QA/Dp13r16tyCslPiXW0fnObBqPqqhEMZSKpY
hVqwV+9/6c9zE7QpDgWq+N1fYDwa45zgACwcWUiic6th3/ki855A349JyvmZx3olRigmXXHI6miJ
7h0hx+ig5eeXbRQHxLk8eovbcmw3pNLH3EPvV8bIhBM5eJTnl5F7v49QoZ3+83P6iLNNIKrM2YhL
0fDalLvdj36F83ufb2i0Y2UA7thUa87lvvNs8UMQrNLHdg7ilhFMMXQSAEdTeF5VeNpINh1Qh01p
WwCf13ujdnAMn46XwShznLVDtP7srwN4quGjXsN2S4D0fU9k9V8T+BJVTTjrAUGfs6onEUkDCHRn
48XN5VvTW9e1eaKLT1SMkJo3CB9QUGRLHTNn1DsGBgEu6GDmNHwHSuk9b5pT3UHr917tHfb3Es4x
RBs37e2+r2k0PPT/qTYU2jSKW4Fek31Gb5sjZ4gsFKq6kGa0xrhCJ/2D6ASg+F062LlzcLjybcjV
+82i9eoaMpIiyaoee1Qkh6hmgNBe1AKuYenrVXQT6xTyH0kMKwnjnajNSaXRoJKWpLG16X6pccwg
wlcjWEgdwjN/WqPcqHMZSkOduUob3d7cv+z80eEFkztVh1NhVexs3tCDy/8j7MVh9zLt94gNsMCN
ETqOabQZWRH99LOJNTswnK9l2lIU2xeFPn2o8Fpp/iObjChyn+RCCgvzAdx1OeBJ12LyuRFw9g3Q
pBKKPRj4/S3355VM4EklgHRW7EtQWDMA+H/uScRNKRcqMhgZdc2TjP4gdt+eo5q8HU/l7Z4YH8RY
p0vpICH/ujYpkmdipLFR2yJZoQPEAzLQG749TpviabR/VK2gCYY5lvJiuzv/kqYcQvVfheI7a952
Zmv0da2k99RSYzbiyPg0mWsPv7etVdslcNEcA6hTvE6ZT1Px6HebVv3+dY5nqxtPW0H8drP+ob10
jJiV72ciXtn31543WmC99FGGYZRqsKv36CYFN3VXw8jCEmFqsJPs2fFUc3PeIUM2fHpeu6OE8Pmv
0Sft3pRfFULoQeBcNGqSJwOdfjIJThAd5mokHKOuDpfXNDtTb0xtugG8gUneiEMmBzd2+w1YARJC
rwarYffzQoYFy/idUei2A/BPoLkGTOj3gIxyHmRhRgZ/0wVROClTvJWJquQQetzrV3HoVnH7/0kY
7JbiDyLD7CTeV9ZVdvIN6lzjb8PyqrHOfcCAZF7oXiTvh1sfDSgHtuktrWOe65IX2mVeKX/4iLvp
w9R3PK5LzaEzby9ws5qyGcnNA4FmPceE74Jxlr05wUH6vO0n3EjTzdy5vnj4NtrR8H0iWM9t+6Yj
pHRcRDZQoWwcgXw3/L/KbEgFb1MUQP/zqAkq56/04h/L8dVenilql9xLQJ66dBzIINYSVc2djDSg
GR23vxva1YLcA9ExYjiQD91ReesNn/DEuMg4xxivbMNGz0UK4IAxqi0T6edtZMY4/XkRq6jBSTlB
gB1b/FEKw6B4Mp3cLv6Qof1up373dbfqKuo/GMpnV4yd6Xp6YyDg6RwNi6SXf+om1jAylkuLmPiA
ZE523bHRte7+TAfySc/f7jLvlHVNaltp7jLApeYOx+mRZ1RWLqkK814n4193RYkAKp/Yrs3FAovI
9ryi2H8aLcAA3Bb8OkPzfjbMsICNtezU0tTr8Dedch0q8ou3c5zC78sU/T5Qw2GU2qlhcpdJo+08
M4taKv/wgIWvg3tUflwAqAfxkSkenKIHfShZBP0dc9WdIrKph437uuKr1wusNCzlrhh8fgTIh12k
UqRxZ8I/yH/uwQFJc3ULvQ5rJNUN6bBHd9uBivN4IvrVuxIAdiVSVJvwIzId2i7gGVtVh4Aaa1vr
+YJWXJ3bfx6zKf0XoNqfDulHQdG7ynEneoVUY7Mc2Hk3yw5iGyKxXk7objVnBdphdIsc4RogZ4VJ
Tk1Ty5kkgISb2qYY6OjRloj43Y+9kGhLrQSGYfqA6d1kWiS4rk2t2J5mOsCRE+SWGZjhjNjel5q6
BQeZNsIHnoANVG+wjynrIJbqmdLKplYnLw/yy1F9/OmZGZPjMLOs2oWkYPH0z2NjYVX0BL74yE0u
JOSsZWsIhDLtfaxlfGKV80i08V26rHRkkJPkqOHts+QWu6bOtPbWsTt2Nz8CTlO708amIQNS1ZwH
QNoeFfCiP6Y/Rbf7OXqIWuTCmECdHvYKf9r9BR6hF2NJDtWPD6v91Xx3s9kmLnk7mzkFN5eG7xce
xoVoPR8ICJI7HIdF5rh4ah0EqtHmrnoSz8IiHdX5yoXGmJVbbIzwtuJIQuACoxuG8AkT6AzmIGiX
dByim60EEn4VAFraoFquPoUAvCWq1vftHEDMPTymo+OFFPcX7h9CxA8v+WLT7599cemvRfKWHqKY
ok6ILYS8AtrZoW7bP3t9NiGc3wvEBF2RZFjEbWQh2fuETV5AWqzhIh7z0y1JnN0vSaOH3NdGUJHp
yIy+xunADdLL+3x75hZuMwJkxp35FSWDddKnv2dK8EcTLs6syP3lMXBZtJdw17VVoW1LyONCY5+Z
JNaE7mAdZ8PEhOPLYpygsnSsYAfzK2AwugvwVDzznIo/odlnYHeeMedWhFHnL1ZITHKzUBfCGKhq
EoL2G0hfleJgERKupSF2wAbIRxZUh/eYjJlIiNHt25GP+hk9o2yg7yufX5t8sWCc6OdG98rkU9qm
Bge1uudSODROowQnJ1ToysxeHXT5J5ZZ4xvIeobSaGsXEFw6VIQOAqMs+NxesmdisuQaYqY98Pkn
K1XISDF5JPDiaUPVVYR3gvmAciEF44vrpgcYOTJjUfHGqoRlEoTIgKPdK2caiS86m2EqF+pNO6xX
Nrzh/dfR3EXQrEbKx3MRgqlMBgxM5BSKjkorJmiAh37jNY69Zh7ZXBSD7XamPB1bS5wyQgIy/tKP
I/2AsRj6rInpGCbcTf103/kYgOPjVKtVTS9Ryy98ssZXYSuODgcKLCtAji5UhIYGrN3mnRaQF+XC
f33gXVyGPmSVEF4ka6dFWT2pJB/CfLJisU8vQGFBHcyAjxEWyPJGnuzyF0DWLTlo8crS01MqFZ5N
IFk++Kow2q/ckMm1xoHOpQnEgTO4nApHqg8MQZpIOIjVHiAxVRgzmdFxrTk3wM4mp2EkxwSQs3f4
TifsABaGHr784InXemd2AmkA1c1NcvDVxS2+Bn+driQ7tT9+8bD6neowhGO3TQ2VmPyP93cw7zAu
N5SM/V6e9movAq7yuzTd1ATrtNonVw02Y6kPQkJOV+4rehjRCEDTYNCY/ggA+RCVPYGf5104+/5J
3siImqMrLRbnf0CF+QaVAU/5vly6NcTE8Nb1BKon2nYKb55alHcH5++dIKKyRHawHXFWZETu1h0A
BXa69KBvzPivc7t5JF4vi6qERuG+uo4a0zjff59XJ8IN0ncGK5D2oz88nhxec0KYYSYL768vKXZL
7B64B9QlZ/z6WJJaQwmQyEN+0KpBZ/WaGZv3g0gp68RHw2Ip6f5NWbE+6yIjaa3zUWqyS0GJdLqV
PSNT9FMroaz3dJ5/USgox8QxBccWnowwFLVdyJsjvz1dc8jB5/nzVu/ddr5Bsg8jzW+p9s+JrorB
Jkm1KBhr6pCV2TorP8hEHF2osRvezTkSEGAVBOYsV6AQ3FJWL8QytaQYqT9EtfxA6YmC/Ip/PjyX
b+bUPZ1ztpuUPI6us5Ob4m9n2M0rkPv2wN0eDHvAEj9mhDX31Swf67JeXR3FpfMi41fonWEi98CS
1FKwI4W80nC1pwomqQVeCLuBwILi5yoyWYOJ3QxM0W4uzUcS0DVawmUf106ldM7OdAxlud4hEe6X
S3zMU0tYo2IMnkqYs+sys7nEUb+eZ9No9xnSXI9mtCahrGDZuQjlG/7rUCBxRMhvG8ksOU5Dxkax
JxktTl8VplVhu45PRjN6L9awki/m1XRMhobVsMKvnPgndzMej4vJx9VbAzToktM2uJVjKNx8Hooy
pqZ9oDSpJT9JKixEk6NxUIyrPmolCIsoMyA2kINCAnXCUjwg24TkO/hreYbkQ6fEjXs+ngnBtdDy
sRVLWuc7BOtFIJ1eFoOdInne5yZBQhpECxWMxGFB47bM2dGhWrWgZOpZ0cuRZ75rvI10mKhNzw5s
23UlM2avX3ip4OIRNPKldcK1iu8fMitfx4X6pfu4kKA+4BqCiLXftB5NlJnu1Ow3CE+r9FIxh6Gi
JJ075EtIKjdISBjXhwp25T1NtgldCKURkEBVTwofyojzxjXcA3YPmX8kBFA4oadHA0Xt4XeTp2T9
dl5L05ahXZ4sIbkzUvTvXJ31+Rl9U5iEuSNmYuwdruVvzkPuCKvZvP+zOaY6ThZ9oRrGMw1fo1Qq
CmM5fe+wol6ehWR5QbvuK3i/AZP3QQ1dXRZuCH6L5LH1GUvrl/YeACn4ryMjt1Rbclb0Vk6/9H60
dz71TF0El8XenYnLr2XkyhiQwySS87bm39opHTZih/eDhknQBXeWKKxpH4ROIY8W89NwXZ11bAZp
5KC1VCiAGky+6YGt0y0BJoUby+NrrF8HjMFpccLgs1/dUy+E6yrnbTkNBzH47pUtTz5Ecjain1Lr
9SdSspFjo1sYb9guZgfe68Xiy8j5vOu/1b+klvWPe1vX/X/OIxNLWSWgTrovG1fDA6/CrJcyIMY+
V1YMIdCCB318sdzViUFZIXbrnEnHjApIV4fLEcHQpMpLCAXh8hcgUdFeuqAvvDpGPUvSQciEm2VO
xyic1OtK0sjfogYKQ2BPfDRXsVng42os/HRtj7yJf/rxF3Lyv8ntgwBtTnq/yq0CjjOR9NP4fCrg
Nhm+LBBvcSpncrQcmJeoDUyy3Ecfsi3ZWVks2GdG5XnsgKVn0m8n43nDgMx94pPD7bSi1LuFRo7x
iquoXFibFupVMXHcztaf+AlXxERvOiZ9VPD5i6FyWxEVYwi9rwRYI7pPsJGk2UgsJSmXcScq08nh
KlMUE587e4dV7Dg4fCopzpdIEdCGxdmM5hKgjI3ONyXcLvs6pbkPc/K5QBYKjL5hn7inwuEqGkOT
DU4KpP4879dPknLcG7WVT2Nsn0TqP9ynn3SYmQnzDzralzzFE3rUL5YqzhkE1xM1J9OB1nUfo5bJ
yAGD4Iv1lveAkYmydGFYujbYNnc2Lrdse1RUOum6OSpjbg+OAJ/+yMfBTP3OMB7BwXoIvk3tn71q
A45errmEtsfEZdHgCxeDEUIsp42KeoaAtriAW4kqOm6MKJlhnGCqvsPELGo4TMRxanQ/h71BmSre
OY0RWz81PTHqZTWi6K0gCwljszVF4zEU7nB03loBzquX6Y8rSx3LGXm1Fkza55WPZRyz0yuAiDeC
k72lRgBOnx6uvWRmVfNBqSYgCwhBBIXPmVKkTAqgY4ee0zP6kxCrBLmlysVJphODvdAnpgFmxoOv
/BYer+Gfl2lxZMsbG7Pj5mNhX54wbTkGPkjlmmTZ2VswbvM9fLVljEz20jVGl9Oh6aepn34sAJQu
LDxReXwv0k+D8etUhyHgJyiZ75SXAFhfWO6APil7kbIdILAbNsxGQbVG+GVe0tw2bsG0/fLU6pj9
AcAag8mmFgRcOUAMoCiMGtLDaJ7SkvThiTp6x7yXuFRKNi5/0tLOv2OgN5lcrEYBC6kr5Kb4tOog
n6jtQMT/SPDFWID2MAh8Ms/JaxeYHSjMk++KRJsOS611llcbBe/SdznOl4EhlAG+KxzYJDLoBwTx
zr40qPpe4NZLjUryvSQwgojDomSuOmZcU69utOUpvcvrr9bUc82scSemUENAZ38fzlqd5uwjglmo
vJBwnvtWo3Nrvit+xy4lN+3vlEyiqz/Z6Q9LqinZ27ns3fF7IRPBIfqV4xlEYUEL5AxGNWBmJHWI
gL55YLr8UkFHtr2n7puVHcWkbisdBhAKOibSqJNpUxkpeGfOXmG9r69wIAwuFAXfDG4AYC4F93xA
EB5xudAyNWef1uIv8Coz8eZNN5WSIBxktcgB5H86x19e2yJuRCLWJG9o7vWusLZDKPz8UaBnqA+Q
pnbE03KQXAQVspRrYTl5Slc1x3wFshQUDWsSzlGi9r8SYDSgF0MYj3Rz4Caj8I8XwvK7BwbOW6Gm
ZukkjsefFsDkpMknEZe391lCHychWVJIswM+DiqwrSq1lm/JEnwBIhym1wjd7j3EdtXrCPbphtqb
GClWeaZrlJVu1lJrox56jek/r3kNRjKkNcRNOFiU+5aEE97iK73U7sIYiKQ8m7HLOtYAIUpLazXA
tixSOsQYNFf9slKJtk7Ssc9cuDbw2OKtGcbhI2ch9E/JRFPYzSIAPnyWM5XLmEemf0Qip7aV0KlD
99jRW/Sauz0rSIPTqxGRMp5sIAcvC+PCnIuzkkL9BNtLmliYtyJEKf6QoxdmlhYF5pknSdKFx3Nh
LhohA3TaWNYFHZTA7+KHpwuCiE+Zj3kpr28qD3AaqBBxftIpz4XYUdZuuC10w4ykqbY5qyDtfH9s
EDNXn8ZdPVhAsSZuvQTKTjWQ8Sndz8ZdKZuI0vsMoLyBMHlRrovnA3hRtTADwut+2bl5KPm6A/v6
6NvsjqCCUSKVq2lyBOxG1WrxA5uS1bBjSqTfVabSqiVpEu7CHAXOVD0lBIu1UK6pwe0tThct0esa
vEczYqbLfLfbItujP2PjH8587PtXdVqQpFKquxSQjfYezRk7t1WRc+AwD1ApSsRSSRmeZ41kZmIj
Qt9l6kegnIZqJJOTSPCFgGhVLZhIqD9b6IoYufTkKsMNRLWUvIVbWNYhQLt41f7pibXs/iMxlhtU
8nVZJ3UuKvHiI3mfqVbkU0EXThbmcD3wMk3SSUoocbFtZIyPtxkCIymU4Y84/3uL6iaaxhUBXhmF
NrBE/SE1hSEFPMJ/aZkwndBXXRHV7/OwjYEbZTp+w0Udd6TXjT1LvPiIxB9srBMsY1DEPs3Plbhw
IJgPlwh2RxlRI9hTJDZxpmNaS8U0JAAN38FeFAjDx13xLv7nlPRXsrLDPshKvL+NDoFqXezFQrM9
f4cdpGGPzi4swcM09cA04qwVGwVKVocBh4VXDTzTqwgKMiojk4GqTWN7vJhwcPY/Vw7Ts1PPEDv2
JEYnlKCTeftm6Uk4coPh28crz3MIi9/Sz+L+8IZ6aO6rzDrUhHFV20WwUdfdzzlmVDCkOz+A02Gx
ZCugrcGZQ35NPYIqjZ8/j32Cwgy5Zg5OnrYem+L+NFt44D0QcNW/vOrAOYUbthQGHiGMepGi1WAK
U3YtX/0HeIzFzSMuEvIyFdjwwzm7d6nfAVAOPluAXeaPBo7NDoAPHmIHeGU3RnKUMs9zHZzSsksG
yRhbS74R8uhAPZpMgG4DUZSflvIw3DIKPrDyMsQ3zNg0pG7CD1lGydC4wEy/gC6+ojvJUKslJKI8
QHKAwQ1LYZZ0IGav5beuh7T9264PVmcJE3HiV9KovAsXGIJY0BmbOhGyT9hJbKJa/XjkFtC9XHK+
MvKwsqXXey9cSuKrgufX5ELDZw7XbEv71fp5G89by1j48oIotAkV0nzWSENUwKgpqAkVLOzHFqb7
gQYlL8Xnz7AU3SmS+/J3dz02KJBpZ4drw+LcqeXetBXkIpp48M9qCS4yzvdvMAr9aNqibjSglanf
kOFrao7GAQwqUCU9tD+aryzOemEoGDCdRimR+B51wEYYkk1Jds9/3tu3E5L0vSxfxoAmZHkiO3D5
wcTxfEh94dykB8Mnne69MueRMeuyJL4PrKPLez6jYJHdIyBFPpBmI9eGXtSCyyu+GX65SIk0Ww6a
wUR5chv7AiBq84GjO4HAe3MnuwcitFKfRqMRPNBlutLhmYuClqS+mt416k4oEt9X9Wiwj2sNy9Fw
gyayoZZhKDTI4xDZJp6yS1W1Lv35rj40tyqp/e6JNtNvDvmJcYMRFGOma8muaTundsWmkHchH7gk
5ZKtjv+E/ax2NRvxlb3MrrnSUKRZ8jzoCy3/2BUl8A2FKpcwoj3qqKOcd59xN1rb2+Cnmbx0SrhG
YkW5JDvoEUGUtZqCTApvG0Qpbz/BvuJqJUfknM5lDLDpT83h0kcAhciV+5lYZNWhffN1g9h6rBy4
ICnQI7nnNtMHLsX0J1hxPGsNY9umBi9o9YKfg29JqjVyRc7x3YbR73Lq+16bNjgKZl+fMQV3UYyw
v5geHv9Hwkjhi9hnBwg4kriPNklEbnl7y+gYyOvc3zNcHzbAlFsaS43CRWhVW5uOuk3V4FKW5clf
PUHi+nHOhbfTA5nN99aorVq3KxzzzgviR12K+gojnRUah3ZMEOzzsHJ6TkpsWp47s/ijVEbJns0h
MvNa/kX/uXBzQmEfI9gz2Cts5sRCMtnltbmXiLlwQ/oQlrZlCM3D/opnaqB+rR2f744ab8iLWO7s
70Ycg459LuC8KNqkcCL1yllcRtxXFerXfFTiCa4QSjA00J/eY3/w2OdUHzAiMAt95xghwy9kTc13
limws/cxDapFXm/BTAhh6af07ss/5SovMFP6Kmv70OWEdkqtLNb5TsAflPUrcoEsch5wgoKUk29E
B93SKgdNXEFZKMoJJ65G7MZBCK804W1fBJC1noIl5+ZVW2SZ7uSXpoPk4qot0pFvcri3mAtnX6jU
ykK49plT1JpHDlWYX7d45xLgRaULUaYegVpw74PjelL/zuGCAzxMvmGaXXG8LBGXSFMk2OYZ6b4m
XRZbjdOGrORaqGyEQW2/haAVf9DnKGf0XcVNtcBHsPsWpETx0Ok1xi65nr5FqyyvG6siOmvGrT2N
lnz+S3bi/CIMHYAGVIMVqYGWbWzdJ7kyCLV79CrKVh4RIrr5GbDwBOvzSZ1OSuQnbnDYSr+kBsoQ
+f9eLeq77zdsYkzSmnWjdolhP5wmdpUkarfmx/ypXKrF3OoyeaAE3V5KVcqY/5bjhy8bh/uMzIP0
h/+GQ/bvmJMDgY5dJYjEDrGPLHHt/tRF5oF7BOiuAGcKYMM+nYT/t2hvSyd9hNK6qDsCbUKSd30j
jcwJVJ3EKqPmhWnUrgM2+jnQw9RjNl3XXOo/8wWO1reHA44qnECwkrujh07Z0tDZ63WLHfuhUubV
WFSu3JbyR0uvfpWszffpEnDK+Zj62hINLzcGED58fjrKlskB8rBl1Zoiom3dbR+JsrkyEJHTdLH3
u83h1C1bm9Msws/TLngzDwoTduh/ij8W7OZtC9Lg51LmtvShG2aKGMvqHlU864IRMJauZgnqwK2p
UqN3t+avne2Sjgu+OxRHhKdK3EX/0GCM19fm4wiupnT5raJb1mh1ze9oiYrsNu193exWtuLc5JH+
vay/Yql1ueK7f/BbS7TjkEXvr3sN5flPDLeG2623qdBB2OweOowDLT2jRZVttv5VcyYtC8OHUo2/
0m4eXPXwpadsmfcl8syip746tXRNbNM/y+AYYzRCBahqo88skEE326HOMi5hT0KQe0W3+k7iL70b
6L4Zi4g4Zt6Ly53WGbVmMEkGGaudGgjsYqCuUe2a4vvBfMyXiV7nJ0Z7V9M9f154UPPFWJ/GuO1g
0xMh3ynjfLvROEOQSrQJqsk5CzODeDh/kI4JSsPkqP459v1iWRH4NMj7jW9+RePZmdRiPPMXr3Gd
/Krj+rvcB1wo8DL8E4lx8qWyYOjHKxOoYGVDsGfkB2Entxw6Sy02RyK5icYATMKW+y5232CbpHyc
etrLhLgEtfmOh284DxN9uXNK9kTammgjixk4m/Aq23yJTq5wjNTx/pfyzKrRBKzsCSwvdCXK464g
TxohM+PplIqKhRaz1SLt4bSfhJf6WJGor6CKC4wx4AccK3ZXE08eTAhJVPqWJdL9AY+pr2mo4XmF
ok0CNpACbDH+rpMFKimU/4wfKtNWIvAv+pWwLI0tG9g+diJRNT0NKLwgV43f/TGtBSe52AvOfztY
CWr4qbG3DJl0H2SMEPCL31lg1g2jV/DFYOJyHCJqgs+kLZbqMyBcqX00NdAxI/QU5NuDaYJ42FuD
kOzLPOThL3dvKGbZCRfBzahV4xOz5P55hf3V9qciMN4e1CSNgxktDzEYmTovtecelyOD8qdP6aXD
tHHGwx/BTKu3V8qyuTwLqTuHEfwmWNreGjK18K5XAoKOJmg5IhQKlr10XQoxtChYPcQ5CpY/j5Tl
DbphCzI9NQK6E5j15qknzf76ZfAc4TuL+eReQOT7w08uPnVdv4pOG+HgvWbfuNK6DGhjf4dzUI6Q
ifXKYgLr+cb8aGbhDITjWMsjB+6kzVUk8fb1Mkfvj3MEFcb3OAW4JsjhEVqCWnUI/RTxzabRjAmq
y6WqV2ZUU70YrisnqNVdoTl/oYXeG6MviA58a0SSOHQoqI635k7v+hEAxdgqUxewRbwYpv40Iqp2
PrMF0M27dAFQtb9HoWPmoQrSyaxAs5N7w565HfTc0dGivl1eoX66wxSv2pzJio5a977oERz2nri8
9+GTIWaKOtZrLFw3Rqiy4xP5ZBIaAGLf+Y6g0oILygLMC6mxRPbpPNJ7W0cA/oVseP7Nn2UXdGiN
hV+ai7l1niHiMYFgOa+nCqzVfwfaectUIeIAWyBxyG8XBIfpDYZ4wnK26FpaD5XB10ZEcaqGcOnS
iUACioYZn6fDUEaulZ36iU30J6bJgkMICr5KmWUM8G/u2QhtWV4lemd4ah8/+1HJ3H3pgxIfSLC1
XD7gRj7BfUbBbPBc13b5IT2hQnetSVEuepVIVU3K4sBEoOZT7GJIiglEIQnxEYZ+oxfHPXMVkv2v
jUiT1LXTPsCMdDHDpDbdEUp73rUgm4Yn9wStbtbGiPWERv7+Xy66dP+WgKx5SSaPFlh+jlOil35V
MOby7+6JcTUDdd8BPL4Ftf6IPwd9WyheSErXdt1dY68VRVIxM/L49yaajMWwtBAVHTCF1w1QnbNh
O9hYqh5UX3Z3E8b9XjdbnNDwmPwXrVEs0YVZSFUxJkxDo0Oj0q8T/o/Nd+0Yk8OnSyor1s28v2Ae
sihgcglJxHe148OHtJuA4TuhF4kIC6iVokhiXquQjGm/YtvizhzW9YyLt8XR2xJ9jv61ACC4/ARN
4TTDLu3h2tHFnOnJBF077XP6mf8nKx4KVodTNYvJL66B8hH0nthaXhZrk8mQ2FVSLE9cBeDwPoCF
9AblglaWPi5rKqoixOw/Vt6vmNTsnd9O3sHbcac50o9hTDya5NGJQwoh3JHlCRC+n2YSs2qrYnHt
GbBIa3/JWe6wHddqDLsnCWWRUACeGDpjMp9Q2B6WjxZlImN4ovnT0hn733HA7l3kts0K6mtDN08M
tb8dCu8OvuKatte0oT4xId3+hely0mvGFSc0nlhaiddgkEsIhGKgY2qB9pJX7o3eR/j/TzbU1rQU
LqMe/rj+GkbL+OkhYZElo2huWXEqUVAkEr+1H514jFUtMNtdcoRkx4r5OHxTg6yxcosgwJ09rsJG
lonIZx1GDGPFbIFyqIdu72+AVPOVYi1hY4wJeecV6WvtjIRnsmlFDpxlUG5djAHQJrvXDZmc6rHf
dyFPjh7e+o1dKV+Pi9RQhsTcGvqrYRlaqqSb0kTF+66E8liUv+RALVsrt1IVRa99a1MSXiLTKkyZ
vF9hQ2KdZ9TJb6wgPD6/4JhXZAAxu3RTk+10xkTFOJWGAtH1ZP9sOu0keDAGBHFQEopyPUpvipFu
aPKl+rax2GTHlVGvd5A/CHpevlIaIWwsyFHckXGhD53XeHMP6eb3IQSSQAcWkFJoahx5mfQW95h2
y4LGstkBXOOmk84jH1bsanUmHKkk8lD/OgKp69Rv3W0UDeVlTemlD+sxMt2IIilASp4H/6/Nbtbr
GxV/U61u4KiGwV8K8SDPXhdMvpJ7j/0cECPbfsSxUefC7vSe4gdOEtn1aUuIYjdtrbuiprSqtRU1
5eGX9DazXXlciKzFDuo+b1E5y0Zb01JEx5yyyoymYfAROfK6zCnT8KvLnZe9zumt7/HvUQfEqLXq
O1IT0ft9yV8QTKRuh06FZWEbNittFqPc4vnoZG1Z624ebCJtDwcZjVZPEhxLxgN+M8gE+CXWF4Kx
CiN8NLXQtP3oIZ73aezd96rnOy5f8JVczfDWsmCYkUe3ZlKRkE0DVue08YzguVoy84agNEgvu+YX
KaGNcfty6hUgIasCFd9QA2OELVdE/5LhePUu5jumbu3u/RST05tTVDesdogsQyL+EaHXSVKMs3r8
qiZohN58Jz+2qSPURtx7S76avbxcARCLEk0Mnjg7Fj5NquU1oRj54UUzg7czIKcUsNfWJEayykHD
F+SKsCQe5RXV1yWmeTgkVJoPpuhON389vcV1HjVm0u+vrOwkZIS5GMEf5go43J5HjFXHAzc1KQeI
VWdhL/xzzEwGsCOOiVuEruGIHaszTfEMBAFacCSB3qNCLhZyop0ANeNSfdEVdTZa/BbuhP3HpiDz
Q1H5d/PNxKZiJvOAKqzbJrWTgBOsTnDWX8/hkkB6Js5SFtyrvV+CJ16k96P5DLDgkBWG8fEQ8CT2
8bkhs6rfyDhjDGd2pTCX3oJuQ76VjQOV9qwumiryGU0X/kLfdJaLxvv39FbcuHdF2W4PHW4oQHRt
vcR5aYaaGHbSqUHYnKKTzyvAuwIjVuOTQncXva7nNr4X9z+qvuMYIL6AL/zusfZtwEh0oIZ9PYb/
UAlj84ghnDwb5PWwJSEWiHZ7KnNcKdU4gUkES/IkbZIsvjray4URgy5X3VqBedbM7EDt8gXeTyaz
8Wur32F9k8zQJ8QZ+EJ4cUn0kYIUCYtLclQP/B59dswAmTjg+1E+t+pyFTM26FJdra8NHlG3FSUI
wL6oUBxj28sGFiK89/Vd+CLojFz5sQlWVMnBK8fnabHsm+z07XVfcgKUz3x6JP40W7VuyrpZBcwB
XwhGfHkr4zDP74BQ+/E6jTuYzuzzZTo/9H1q7gY8WzQeV2SncM2j60FPnLSmLEkD6A4/io64KFlm
UJZdrMaNyam6f+2zRkoQIU45m/2qQk3Dbf+NyfsjS+rBCRxK8WZoUXiGdREZ6Dv+VOTt2JIX1DAz
DZa8LKFbcKGYbbGjcq+grJ1TDvxxIo7RKugcGxCiySCHRjIarIK9M4zyHmz/EX0utrxjToQUz6kI
uAfdTQTj8axO3h46byjMXuLULB9XxZZcWYTm7bMYjPTGTZHm7CriTy05d6gAhB20JNTkKw0ZdUkd
kBvEIci9z2EFU9snLnsvcdOU7RCVG2J346c/BnDdwtNzCDWwD4j3lH1Ce6cu4Hx0G2C0FZsfwToy
vs8BEADwSftaCXnbN5TC0yfNh6vXUqF0cSCp1Wf+ug8hh+J33kd/TecTeeztGuC/v3ela9Tdmn4A
awAxdIbeaqiB3k7L684NdmDm17DgWdTeF/9XDm8tBfNxBKtdivSQOjrBMSuGTvRN7JB561fABWre
mQrJvXVXNrQfmWeYbL4DaAIwu1tET1gkVcLe8Ht7KYpYRX/TE6fL73JupbCAGr7hYJNPwzx+5LPh
KRej3MHiylf/Bf+O0U8cXi/NKKsOlR5HO+v6CjGNorlJbEN+WERCddWj3p+ohFRwW7HbdBuNSOuo
7d8eWAPau5Fo3YSHiS0TVK4TL8mpaf4/SEbVm3Py1VvqPC10YxHVsiiaVdWQVSj3H6NS4e/yU4OE
DSpLMGwrPWrmHT1MFnPpI+hv0aJGcyFqx8Nfkl/AIbfC7i2QaV11dfOOhEYtzVKdmCWLbtUZ+uYA
j8elPpbFYJfYk9Qn7h4aJ9XVeMKZEjw7Oi/sld7JGg1GleoUdtbCzE1sReYhdS0zegNJRbSJYrNA
tZHhsFMzVFoBBqbpy9qUOgYYWOzxmbuVCZ2Pga/F7ot1dLOP+XctdIJ5KDttC3kY5sqa29MsUz9m
wNwy8p9inycuPd4B2CbttTytnktXGCYJq/nsIxipsdt01nqgG5Vn8QWbCNJ6YVSsCGngrxpIOsqV
yQ6MAD2s6+JPJScMgzPaH+RARs1QjzPINDufvDVyvyjrfQUTO01+uTZvqn9gR59nKkfm7EWk6+13
LfmIR6gw3qkYgKKwBy2MC9RltsC5Wbl1LAlgjvnn/cHpeF599eLACRJo5dsmG/TWju5zdGXVPdpz
agWzzVvlH2k5if1+MAiPraIWEJbAuU7vOS5HqJJeZ/DGL7OapCdg0UfuznnrqEwl7jFrKqguXeG7
RDApd501YSIX+RbG9W5K0sLhTvykI4bxzhsX5FeO5l0LF0K+o/VfNGaM9k3QSPWwem9f7PhJDQzV
RBeIy4J8qVqvHscTmRYoALvqxwtJPDPkxeyTDVZOJV3DLKNhXo8wlfIpXBaf0jouuRCvMpTSe8EB
XJKMCcikPA8ke9J9t9qXxq9Q1LKqyUPj9aB6dewsJZR4gCm89MOLeK6B98rygqRX6eN1vfLU7sgL
Opbn/KMi1G/CKzn6caQ1YNINqhUFXZ+oBuMg7LUIVaJReTUnJEk4rmyaGxc40zDXwRYFXcUfQwLf
CWHoOiw+AVMG+x5bINW7U+z5Xubjph1LZ88y72qwuNHAx1UIgzVAgC4QPtqJz9MXzW2vgoB4/8zO
JhD9yi1EZQLRWCh21rRnk3fmYYaVp+SigZdfyaESTaMDRz9QChz258zHca7WulXJEdYqkDr+kT+k
4KIvBopeQEofebk74VQepK9jNE6rZMHD9/U5TpzICTxiDoyDeoiA3ao1R9XWOiGZnLcBx3Ddo2Ci
sL+p9LlxM6tyVQxWBEs4OqpO+HSsIBFoKGCc7FXxJ7AH1WVycLjCjKOFbb4ZDTMI4M2KOlsIUVGl
ivm20HjMbUSCQu7G6DOYZwCib0BeojYGd+DE58JxTa7wA+jMR+WX1m1gVv3ruqzDkDE7SFKVn30z
c4KlRMcUpRTIXScFmM8WjPGqf0Cfx45onj7rFW/RQRt8u3A7u/oB/BYZUCE+R7vOuMalNumaRafE
JorUUSZWFkWXNSJUeo15SHSpK2DqjETY6Kq4eyBVOkhXqjAWNnP33QP1eTy1HtE12yQaamdRWCJs
7+LLAZV2Rh6kld/2mvXWZ9Dj6Kdd9SlrfFa7XxxZzTjrZz2la5mfeCT7SzyTXcYX0MAWZPn1K2sk
ct4QNYMJLPdbjdIA++ZIBEwCotmDftsEiBiF7hrMcumfhNUxbqkVQz7KiRg3AbiFpFXd7zvE7bC9
JLQ5eGyobP1a/aZ/VjqsTTGVBhSi3m5Zv1h9O3rtOACrHPtW78ICTWK7iIbORvAvJAY/pHri2bo7
yXzb0P1hbZZAtdhcYZjL1dhyhEJmSeu2/I5fKTzKlXSj+HgsGWvUZnGdAUmz0rmgFHuCaHB3MsC5
LufHTxBFow57lChgrRZM66aAPyNghwoHwiHZch+qkADhJ8K/Nvy4mCrcjAmZQdYUxhb4ELfd8hO7
2xuR/gjVfAiekg+tgLZK7kJnaz94x79gMCe2ceEdWhC7HL93KSBV/Y5YjHXwnbilaI/7+e3CW5xo
pMjJ0nRlcmEf9TtLLiQVOdUaKCCufdd/ObxQll97sZBx6Fx6CddMJEStuozhdwdqaPBLQmBcAbq0
tFultDli9J1P4T+OatZZyc7LfwjCDXn5z7c67XlLXf6+c9dxcVk26pfBmnPROO/DUlYT3qzMWLJb
Z5v3qzsd9ZgDGwY6UiNLTBls3XwfnZjclN+QRlnQf+F95PnhiXjLrvJBpNXwj9LfhRr4vHY7ZD90
a1kBK59uc3X6La728OBGzUEVxqaA7ztYKP5N5XtK7bVAzeJaD3E4c/jt9+pa5/+6IWL9tkQcY/wt
QjcpxzTyCVeB2KWsfCEyuJfbbPm5KciLHIRoKZPavW7GfRykV75GJg5BJPTFHWKiMAWN7lrXRG7w
kIcyqySawwlJZ7XAS8/c1pNlZPIvt04AJG6966qqfJqtCmZqx514FeSFqCgTUC3uBlM4aVcqjwdR
qwxabDO7VpaTdZL/tXAID7ZryJg4SSHVOcge89q1z1Fw6e4utYg3kgUrCDOlohydR42geJ3yEhzD
j0+HbORJNhea0BJTuSqYq7HqNj+hMpQty8K2oWXN3mRSc3W+M4D7Gi7Efg6A2GkrZAO2IBEx0t94
6SYj3VNiRQSUEKYZAXJ0CusfUpze+pi2vPgag4EB5QbW7XdCyt30BcEqbQ4xde1Cmiy7Jiul91yA
E0fNA6mqIedplBLXvOpx4e96LcqqSd17ZzmRyi2j/cy6uv4r7ydRbISRzJuyXIeDtf+2hJXpZE5k
NkRc7a3ZOtEMAG5fh13tSXuC2xb3CcLi5tqrZae41UBEVXManPSezXp43oQ5ylBd427uCeRUbj/3
CviOVOjmVl/+uVM990goBtzJ1CdjmYmxb5MF9fC+5YcreOUHn2gBt+AiuSphBZrzGm95HJr4mlfn
/1/dXmtLl9IQr/IPrN6YDU6vEGptjRvZ30KTrt/zH5+s7d3u8V6tJDVrxSjDwkZBdlYLpdf0Ihox
zIQkr+JjWz71BElLsCccQBrnDYhCSRHbbtKO2o/EhH2OrBsH1zSDoaIvPK7FnE+l7CzP1FO7Oyww
fJjJH7DFowrr+XMX4u8mvVJGwC+/J3PDI9Iqw+cHAj5zkJIcG4yMrsCOWvk9fFEBFrKONHNKpUpm
WSunXUk7w7sI9hgxnfzI6o7wuEK+wOCUN+nWyHOKy3TVHQrsSlV5zSlnv4PpKKEILCKP55+J5dH0
73huTc+H/su8whMgNjT11RaNRvLvnjJJQcUhVKgLqgsY+Dn+x71foyabuQcYWYZvvINIl4Mocs8u
8aNCPXp0nK3OxdS7fIt0AMsVLpTSXstXgHk3H32Tt329G8+ZQhRUqdSt5JFaSw0QL7nWxBjkHF3V
FS/wHFKlysZ8WAM7XYiQJE2xrYxKWZgd6GXcCQpIJ+GCNFeXzsTRq8PsH5vvsuwKNhaRL4ctpRSX
4BEwLTVdv12ijWtM6u8xz86cg4pFZ5H+c/nihC5dABmVl8qFph4EsiHpHQ76SoyuUHzsNkCjBfBV
iyvJVeJdwTQguDMU3EnhNda0NfjU8VYg9YY/S5yNAhUNOO9664S47St7BCTjltk6ZEnGHpW5vQow
INb8P1w/nh02zQY9I18QLq7jEXlLfrAKeySRimanXb/GdDcf4krmjR5ge2Q4n+DRmGgznbqXZUZs
8YfWFi7wFx104jB2Xycb8j2jUSA3R6yHWGyWkBIIuHFqO+wZCxtsCGdQj1xCNbsWW38EepZKGV+L
9qT/PQwe0NrAe+/UCOV4qCVICYEPdiZXQe8MHtCyHhus77jWDBwrr9KJceayrRVq88Z6BDFXAqhz
Te/7lLACmUAq3m33k+Xy2LmktB3kOxsFSOOHxMa9khQz1h5FZHYUkM2wUPk6e99BDbuW2dRimWha
tkeGzf5tRlZvuIcrfzvSvlckojG5o8sCn2oiIODCBEZ0ZfJCQWD1svaO4zqEuTOw0zF4uwMgUJAz
DPhA9TkKBrfrpAmIdvlpi2LrFoaONlPAJG1CB9dbbePvru33oR3Osq6YpBKmr4pAG3xqxVemodAL
xWdk62vWz07JTCiQ/Wih1BczNvqwZxVJWDpEyW7da8fhKiBSd/+o19hTJii+I08voUXxpyIoLYy+
j5+zdVsAmlgM+g9ZwfaevDhNHNsnU7s0KBHArc257owwz3Cj+luQ+Z9RYsRI1Ydy8IDKQ9y73yUv
9IGwyV2sMAI3O57Zb0q7ShTHeuoKaFqdtWRxlDtcjRS7oixbty/6cjjSTUuqyVDZCxLB5oos4cZq
6mjiVHbh94N2H4m1Bjnq8QaJEzIuFXbH4asuNj8X7DiAnBOfLHYp4KpGZ4DS9HuBsUkCOTUFYHGL
+knTsyEAu3cgxRrub/S7FMkYjLxXdAbWVF3/zUBN6hh2AohqnW8H6+JEdsuYRIQmh/gQcW5hrafC
LP3kccVxBkF4iXY/j39msZoDIJ9pRL25wFwbwkrusZnSbGfBRVooTTxkM6y6O5+36OWtALdTrOZc
e231HCwuSQszDjOQj+bq8xgvJhErP5fRCT9YdF8DkKBK5YEl+2CrxamvyUu7do1ywnGSX2rRCUHE
AYhNKGUaMS3BKffON/dK6umkUiXAG57xqMGw6b7xUe97ZPknXgsV8sIUHQlmS/ORFwbtMADMMhxj
yypckhrwLvywrEl71G+Q4Sh5dT8uEt7ciagpgV7dqjn270PCrw4rgOGH15EL7jYNI59bfPd/MWu8
V0AQ2L7HQZxvGJ0yvYAdlLnjJYAaNl/6ZF5sq862LiC3zyBg2D5xuDdbdJO/W+WD3a7MfOn2Hz01
wRvlI+pvNvDul1oXLWYApmovqiFVqhNItkulTzukUhikYgP9ufRM1R2b+8bYPvvquVCY4gqbmcfJ
QIrJWcWbdLBMOpQYVflvdJypG2H5u12cZ3CYhRdEiqGeE5rS0zcXhy6zJZlmGpYXVU/WmJ94VWRw
p+J3izADgidub+PVeMsxIi/fHYhcboYEnEDzUgGZ5JQ/D4KroAhAk8PX8M7zHbSoZyF5QFHeQStO
o+2QIkT1nl8kFWnk3mW/RhxB/JCeFPOs5HwPQ8HvEdKwhbwTm7lqf8Om8C4iPMRO7fbJF7UWZVLb
lr54z+ATc/tNOkidZChjLfOoetZ5qdcJ9cpOP8kD6SetJ7d7AOwu8G4hu0mehDhqEnhoWzKIp/T5
00EBTqOZyhchDQpPlsS8THPUZHT45pCA57SSBKQjhvY0uSiNwSh3TI+4Fcq1V62RR2VufaOvxTTt
eTwE6AQLJsg4ohlvTmdQjtWq8AQk+7ACYWeN4pVlZOCsoXAhK6Ia/WX9jSUliofxXN+THhrVeF7z
sjKGozCiyTRaYEMLBt7Uxas795sSEXrxzVGEyUC2ztkTkrR7m1e8/A0iWBH9ZAZ7wj/FR40q9+FO
7GHly80W5lDUIdrkM8XyUSu1+84/p+FPFZVcSwL1Or59V8vWi49hE3eYttSLz/wKcgoeFp5MEVr7
QaXvOZzvve/y6oAmhHBSPLPH0DLtYNSv6YFUd0iy4XM8Dvl8HTPNsyQbOSV2eMOOXPZ2EMETgsuk
kB3CIrewcl66B7MBbYTylzMTetnn0pFXs2MmXjpZeeVT1opImKNnCm5IxuGi1gruvd4U6QJq7uhy
03Lh8tEdQY+JhbS8WOOFhH/YU5nFzAQFJJ40tj28OpnPz2/zJlEorhSnVd8zxxxbAgXX95mww7sL
56cB3+KkX719Gig060oR0Yj5LkFVx7eXVXyqJX1DtE7soiLhYEnLF3iTOGsBScHME/con57gU/C2
PlitZwQH/ev8N/pMdFaeSlouk4Zcpswj4baWTf3qLOKsi7kTWyRE5W8X8F9SECbZjJSRhbeelRda
kmq3ren6nRwjpgnUkMnt/5/iZ7YoTuFZnzBb1w9YZPKFk4ByFSYZl8G+BiC+ctdxpP6MZTnfQIZW
plmA/pB+sysUWxZOq6MqsK5jEOmQy5PDQ+fOECL7+On4p87CGseNnS4HHWQyXB6R5l7cGtFQuKgv
5gxRImAM/iyETNESeih34CihoRn/jyuFe1jfMl6vzzHanxlPSONgsVtdgDIBh4uYKdJDKmhb6GuV
y860zS7jpcrrff2mvFD+p5dsIPQG8+ZvWARIEkPPLMpiPXVsaJ5OneyvtjVd6s17/PYJ41qe3Ziy
v3KLoSmMDkFuuHIz2oB253yt/yM5hVhP0o7tEzwg0b7cO2efcAi4PTDjOdOBF6WP6Tr8fJIa/Lkx
+9I3/1D2s2RnLbCU231qzDKWycRU7pLk9clcUYRoalcjErICNuVsQpbCQ9joDjXWr1CX7+rrX7wL
9xT68B3PQjYLSowBZpLzlJvrmTBXMOeVQ+ryfXCvQmYYQPdf0T4oqcAlgi/Zi6cUgriCqQ/ZCqXL
0SUYN6U9uEW8Y3LkDd/9EJsbigmHOjPWkcCEnsa1wT/kOleO+8asZ+rcPrzUXJgDtSWg0II7ZOgj
+FbKxLlr3iPhd0qTTyo/hOx02mboUj/CFnIqiqq7dlfd8N0uCV+lLfhJQWwkxzkG6lUB8NyA7kug
b/HxxJgyUbt4oUlMdXS9x1/0GWBqNXeyCdJ3DIYqDtTFM6ogPnKVOewAKqyiliGCvUhhG9Yit0Ji
yI6GtzujbsNvyBrFSigy//67upoLAzMIkZq2nRR5FJ5XNTaQ8qAZXl7/aLYjYD4Gy/9KLktcVZvn
k07VrhGwpPLJcrCJPchl/ChiuwiTC8C551lNRwYT2hG2PmkbuIluZsDBr9epC2mFIxiir0FQPNPc
GNK+A7fpZuqSG4PhaubIqsHvBmLId+vlgK5v2bITh5gkenZUdTTcOduk4ocvRqtjDR5O9MGDVlmR
h/ENGnF2/h/Nuev4FZqGcEq29EdGsm4ZeJfqlztcALPW3jXh2AaeNw35TfE50tBFr9eStPUPZrc7
jaiddvfa1WtnMgbGA/1uAwpSoZtNh3+n7F56wtUdI4DIY1BcHsN0ZNfTgZaTzkVecer5+lQ95LgS
yb6pSK/JasfSj+yRy24DkF/mTLBaheAt+UVvVIenSV9ngi71iXWam1pROtOqm7L92SSFgQ56klQQ
E/zqPEBhy4VYBhRBcFArbU8VtouWo34HKZ1Zo8EKfDnn90u0BZEQby6M3UIJ7L3hVe3idmDCdhpx
PIOhy7Jbm3EC5l8iZE+O09P8nbQCediPWkouU36H5k6C4u5MbD/b/G1rhB78sZh4U2GuuAn/ni66
Z0++1wgLXDkkpBPYB6axApKXiyFAs6n9OSbJNrr4Z3+UhXBBu4fOzZ0IjJwHJFcF6o66pFxq0ae+
NfyHcpjPbVGJ/K+X9wvjPxvZXVqbGFEo1wfokR3SSryFFV1Bpb9qQNB1FwphlYhcM5gyzr5Luxj8
pwdQjMiGum9IsuHZVXQSmMdGvNROiy1kpjKubiBQ1W/p15C2VSpI6tJDjUNwF61aeXcJiSBzcYzP
TJTZkIuZ7G5f5harS3m+aX9GC3Kbs2MIjSt6a1YQ/rNt2wY96IYpkFVy6Bjo4NUjjJBUFvl4Z4i/
fVDvwsIPfoCEStseeNulX8GFOWD7jVLw1AGR09fmhx/ntcw6A1tD17tto9J6WcHacgMYTKDb6o98
6Bc+rDMxZI/MwYaY5wrqQVneucPloirFW1a64DPvjoN6AeA8PbD3V0jcxsHmRS0H6Ciuwup1T3nX
Lf4KOJgnWidZuBaWj0b7dj3cDIkgd6DwKN0yar7BfrQIfA3fOk69U9j+/VI9LvV9mWA78qrcBE+c
+gboDZCYI7GdBugJ98eNappJDxs2G60eA4T/8Q6pBcc8/6dcz54LomIxCF1qok/qRfdxfkdqow6q
fwBgSO8l6YiRpwN7sDW+as1Th+OBkHst2HaGJ2S8MoYOQ5hs4llQ0SzjQcq8uGAXcsH03HwTvktd
cXLYb7/VwNocmMzsg/LpzijPmJE3iwp0S6ZOZpK1A03SDL4lahOfrIjvw9jfFbAq+gC7YNVy8/VD
tuXjeEWXQmsgZKRsMAlPRREdnNXPOwS1zzQzv7u8O97Jev3mGA017ZA2wgdmK7FCPTjr6FMZHmMU
ikXo4SLjUcsXTev7Iy+LXsNsc9FVp73wVpWbRya13ydWBu9SuiWf+yiuBR3Rr4wbyPuc6d0EN3YW
v1xqzHCVT9thDTFVy/Fmu6EDBzw3Al3fwS4drDhzUmOQnlB/G68uWbXh8BoCnLGxZ/LX/Wfr3oDk
OppsG7QGk8T3IIEG0lhLL1CfuZPpkbt1UaIHeZV/4cp7XyJtzP2a+2ojRKUGod6saJOyHWSbSzDO
8scGfFj81NIJ5mKPykgeB6lN1iem5ZOz07zuI9Gd1WzQ3bYbR4LmvmFJXbKxpLM1M91W+GT+2A/2
922RPEjDCUstadGAKqtQFptc1w29gd1F3/25cRQ7M+fn7sa6SC/oqwFUCzjse2AWoNX/fw4bzTYq
PP8ID04hvK3eekhzJ+dJ6FrJw4XqwysCUBEApa7C6A3Li1XyKYK8JLkPnEqx7wyibHZEuGGp+EGV
2CZ8wlb9rSNtMqDov8pvUISUgSwFIPtLrmfANZTpO0VkEOMcOJQyfdY1LzpXLeH3n4nH18nVfXSf
p0BgPLN9Ca6A6YzEMRRa/b2F+6quyl7R4jIjqVhjD+vsclLu7wrmwb8NHu7wQwYQ++v61MFEv+MS
FkJTQQbyZZFLfoZnllIKLy0Q41LO0eRuzIgyU0S0LILEODbvu+SNBMhieD5pImY5/xo4IeURHWDO
Pb2bYdVvOhcaMjNqSjguG+RZv4baxTMzAiYCxFC4VGGcJ53U2u/hWE+8+MHV4QWQmhetPMHbao2T
+ecNu+umTBJW0+92Ikox8vMPV2T/h0liw4t7ugB4lpeSESW6Mm1EkWo77oGGhG/uVk66RNzCJCB/
4nO45uVB6OXLQZCI1J5JuOV7lf9LINhP3BKRand+Sb49JwzJcb+JGNh4HTESdzeRsoJZ0cPdGyY1
cA3cbd3aWoW7VkdCgCTWaiNLLGPoF5DW9k8R7T+5tFTzketzPAtPfQVh8uKkuwaDmzTnRDvVsMmf
qZHDzE51/00VJbM/wzOjqAGuqZl7GIG5qhe2vewJxqPQZa3RHjkFvB6x/qYueKu+ZwIshg442MaR
H92EDqMpUMWqywqWcDngYD6n/oWIuPP0lKhYVY3256vK9lpyQtWYmx3MMznRGG2HXF62aoqyWg2g
7+SH+cv4cl+CsAPiZFBpg5vbkhZTYD+mJR0f9c6zHsfijWjyFzj1bSF6b+eMueUvIMeR1HJlJtgY
1/pmIIIqmHPNR9UjJJuF/9aCVNqjH4UHdDIk8Aiu5gVv+1kUlW2dMKRuTcS4MQ7blan0DU/X4ZVT
+8se1uX1iibgDClSzfq2CPv2wZxUEd94GPxc2GfaWzB/pEF5rz3ugNAeZWoQc3s/pMf2hwfFmxph
AAsDNtEShdcWPdYwZ0FJe91HInijD3ZBiO3QoCctIU95i52O+fryYNCjPnecs0m84cW/yuiemeH/
ulAacznUnHmZWZj+h7f4S4qrbP9fgwouy8FlIENuU8bIGYklulcEZynXCi+Dvq75Aolz2aT2e55W
rD+nJ29XzHUME/ttHHmV4mI7zNU/yYRxpW6esQQQU4Ilm02I9An54rJ2GGCbLGp7rOAR23um/OoK
HkwEZtqJsiAgY+MNFci7Hn/WwARtdYBJnbduz43wzbnh1bwIF4ZK57KsabMEYVrxQPGNP2lpIdt9
cVg1HhZuTEE431ooQnHX0epuWWSyMawlfE46EpflNprUuEAr3nHatN+Ac1TLD/nRXHxJb/hzYLNd
B4VHy9hymx0H+G+1dzI/YJ8HD4RWzNlOjW6Zm0BAs4JcHJao67trKuCMUpK4V6sisD39Xi4Ybntf
PAjCvXs4vw8nMbaBLfWPV5t3rixztvYc/BisLI6i0X+qtl61AxwbnAOoxP/JKsOhgtWTeWQQRnrk
8KV19ugENd8GiYE2rytjLxjFUS9X8tFctZul74q1XJJ7g4QuFw3Foll/mv6OWZAYx4GmkpU6oRyD
OOmq7O9sstYve4U8HbCc7oZ3IvRLPeIVoMupJEKVzlkU0SFsa5jehhyoMBvWPPXllmfG9WQIJFS3
PmOZD3ki+jhbqkC1pgunOWhc64QlLiXst9ZH8/wsM/G7JWiNJEmgMPGBG0uqklhO/ZEm+9Mp6JXp
lVkslC3AB3lJJhmYHs0E06vDltL45FCDPzB27UqwQRsNXZR3TqfyseHbT4Ciw7SV93luEjoQXsZF
ruPtBpNdvcdTazHhIUw3mZCnIalA0s9kCGif7m2uJ/RjMqrKEK0PMvGyNuIrUgMmfSQCe7cjvpeX
ojxoBBDAAQBa2yeosOl59FXPhED7/TrpS3CW8OsjxA4gS3IlPU3I1mxJs/i6BHb5Rbx2l/otM6+E
hdq7ds501O4XOOOQDTlLWh/g76jEPyj38qHav+HZKrVdG6d2twoMvShCx3R7REAtrUILF59JtAYY
zIwKNZUsE76Aoem3WYubWSkP7ADJnrZ8BEnuS4355gMIPsC//Te9LL+hBxSe6IYznTCi94ftaijI
y5msmLE35VZrMxdgYX6m7yDSz8zGThUN4XyPcRBFLhBmqWyx0KRawNdQTFF/Iml2mos2F1FG8cgz
0drtze2+0Gg+SOEPsc2RBAog3ogbbYl//mdIY6S50+QmTlZZqFgXc8rPqtlTPv9QTcBa+lMKr0lz
4YS/my9EXrCaDKC5D0mgLBnf5Wb24Kl838EivM+Q9pKMdzAVREvzGGZGirrcpqVPHPx4+qmp0l+I
MixhCxgiHg93LSLF6XXeP/J8Bu6LNzxOyd/hfBDj41KUcPN9ZKit8mXv12S4y76PqchhvKMRGIVg
BLVZFft42TBC5MNW8VWgLRZJw0IfrO+hdYR7TwW/lzJfYCbq6C0AX7Rn6u/znZb0Wz11q6XmR4v+
uFaxkHN+G3mthrNM7QsOUdGfGaOFdc0V9o49zAF61lPUIlva5q2AKC2TTY9ezGslMPNbWteAIBpf
D4mLrOWc2rTEJhqVki7B3ZdeKIv/MEd8aqUtz8pKfVpEIdqROVaCckBnsnPBldGeSAagOBUsizVA
CVlqEAl4gE1u6ZcTH4qekZQ5FxydI+kFdp+iyzZZxbdUrXZ4AY+lv7Gu3yxBinp0tw6w+ZADXjXA
HiDjsG8zIZItgKZlU2TvUdWxqJNYjquEIfLUqbbvzZqO+3CKUUy9ImzjxWCjM++kCt9vyycFfBuK
9DMmLVb+kEHiFC3TbsnXUfH+e/bSYNztjWk0+Pqg0czg3xEKb8zUutEpmF9kGkJiS+EcrjbG0SVp
CrH+AuDQV+YazP+tI6RjTFd26A6Xwo69o7VCbKN0P/e7kOegjLGgZr3Pecv52u/ZN6/FOPXmC1IK
4XhgGlo8mkoWk4ziJtsZKUG77/0oVgBbohvXIVGek3Ip4z3znd9AeWhQQ5aLfFuSK8ek8DIdqeTg
sawJk4/ch1I5Tg/kW+st3gVyYVPgErIgoafr15nex2ySXsEQvG9boODuIqOv0DDshjyo0rLj0YiM
Vi5r0xzA492cHIHPZJh/X14c91YsjhjLU/00sLwhRKvFPzrMHenH+tLEqifTzj0oh8YsxvNSekXB
3/XN3nxM1lHcLIV6e2FKHaO3ULqXBJpb75GrapE65F6sBO50QyWp+cx7Kr/mYqMX3vSi5tDk9bEE
1JI8FbYaU52kX1XhAvY293S0d9wSC74BpPi4d7uXsfC8bU3ScgyXsxx5+SAa8AXDdfXDL9+48DTU
youEAmLrYtKDIYES4tX50XKvsgEq6KU/PbI5IIdWAhYkuh4e7sTizKbAYJds56zfHtVpdq/3T4a4
qNcYB3yBmZyEhAc6QUs81ZpfD1OOy/8DEdNQ9X59Rub97tTZywYkxq33fWmWFvo7KLwNOr9cBaEu
YPihY+PIuJeMD2EXS5RqCuHRhkZQTt7CTMkzmpZxGU7AMucteL3WYMwLarmFvhixMOZLH8QYqQlD
eLklzDBV0uCWEFkU2tTcE5NQMbEFECfFQwitiimjprk7Ne1RgJe0t/WU4/D11os9OTSUqqC0K4H6
wKVp1sKGcPw2uJRYl1hTo9XNnhCCJm7MWgM5fLA2kKCr9We1Xc8mknsYVSzOsAt+0xTMAsmaVq+x
zUyj8VnUyk2f9Cyp8fpk0dKDUzFzJA7XOvWLm+SCJZa/YjEhFkr5npOg6IpBcpEOgPWPhB63OAMA
Ko4UvcR0OevduqOobW78cJpuqeuf6JkkYfH/ONOcUh+5c7oPpfbZPEi2/imc9kIAA7c34BxDwpeI
9DPV4z/phtlzMgMGhMZHMGf30eZTMj+o9shmCuXUYlcleGx+k5rLBRuSBRBzin0Scc3WhiQg1xfr
sC7JQ5HdfmVvIL+HKH8R+D910vkW0X5ikGwtzDK4x4lowsMzil7n/hQ7hfVv4M/M7lhJqttrquAI
B1C/jght/mH3zkw+xQtGqw4Zd6N+MmQfQ17Fs4w+GOxSoDxsEuv5pnXJIKZQTzlrbhEPyeF8Om3L
NNBbktGGnVwd7lWpLv270mFr+4g4trHPC6f7mggJ3NWPbIq5yr/PGalQYtv9j+dsdZMk4YgZK05s
q01m9ZY9Ibex6u2Witr7dv3ISTnnJZYaXA6UdqNGyfaE04RiX3ga5dcNc1OmaMDAf92vK5NrPs9a
ZJ8OHtAY/mNys4hUSR1a7ebWvoUnJopBd3xboFEseTtaiKoW0s7dFZNzNzA2q3gDJPi9cK5wOaNl
lmXNDFv6OWAYSFUivOKOTUjR64HLR+0DZHFjtWXMeeJGUGxO29Im076jh9vglvA+0tRElALKXsFs
iLYhiWmUfTNuyRbukKzirD8M6M6ijFC+NPUcvVEgxgVEGpVjF5iJCYPGClhyQT0z52En3CwyaeQ5
Nw7mwPjy42NFEymfVispzDRvmrIAoWdl3J9wzwYuDezjs1+v0iCbt45f7XaQsIWdjIFaq+wIQwRq
0ibly/dZC8tqRkWhhxKcaUBWvT08im4VcSR/3mAkNBIUfmycPkROyUSvrZgfshgWMvjTU7EkwdHA
VAwJD96K+okxf2HfhQVi/sJ7FdIawjHhoo6VNjAR16d6uXz1KA6UjQuUrvQ6Y1LWjJlY193mMbbB
WYRQjjY2Posr0WZf/R1k1BvuVjTetQZLrWqgZ8Z3IIO6JdLo5hAlABKmJHe0O4X7uERtr0TBMq/2
PW7mgjmK3K0/flCeDq1cj/BqAUGMt+TL6prXpGdMeqWi/jGlGwfzlMEjc87kkun6zKRB9Z6LNhxa
a0Wjh+hSuQ2arYxrX2b80twGwWzHSmH/DMRkVu4YnsHhsXKZGKpImGroEcsUqw5gsZOD6nBifSQR
Y11Gh0mDbjHE7xBKIlscRO9RjGLgheemkGVMjaeEXWed5aXN54/rMwUqF3AMlhZhXkCW8HBu2NdM
1A8mZy5UtVU9PivGFoOR1VsiR7s6t2eOU7SkHO9Q7AiBWKcq1KQRjfncvdxjsgoy5LU/VArYJCEE
NahOPHkpuTAHerTZ6vb6HG3BLDC0Mun1VQ1q1fpCrRJ6T0an/8s3E4tcwUZbdWZ5e1l00hwh+N8w
NKwDHGdNdv0FibrhJN7DUayxKTIbqZ8sSG9sb3x36WviD22iCsKRA5iu6m95HdUMamz0Ud2KrfWP
s7H7xbiPOkYVFZMoDIYvtmQY/pFz6JVVvsn5J5GT0XdNN07ZgnIE18a7W5eBhiwPtpfB4MDq5j8/
2vUREm98xA9bXPGIFUpx1ykuem9RFujACKvPglmdVhTcEm7iK8LabkseSbbwzlf6PMzyFwlLqn5F
LoQ7dEZANLntMAAdap0P1lVqOwjeObLFjrYmnD0D6dpyDGBfUlT5vAuR1imEdSwoKhkIxvbYnXdS
5l30r3p4b04Z039M8y57AINMNPcCabCzxyf1648ngw36Kyo6tw9axVjbIpQbq6emx8STRgR8bWFG
maeABFUbJPBkNKrPkT6xZjNCO2PqL228aU4Yp/4k7mgHqLcBbYrSbc9DpHrz0eVeuTsTAv5SHzRc
HrZvBy+hEwm3Ignec5T9qgDnNPo0p8bQgEkgRIziLJJHMpW5t+EuhH5AHqFiVRgTWM338qgb3DTs
e2ybi4wrdL1Yv8vf6dSWB3H3HHxpLFPucwcYoFUDlExvjVSr7B+AT9lFwXl8GAGqYN+ULflpgXfZ
yZU1mrh5StL6Bh5B5RCVLVGY83Zz1lBMaGkHoMZjkXy3DVt/ksn/L42+ggmljXLAVTh/P96IB9Qp
J4J0vbbQzdbeG46kXp54u7d8FuTlQWbf/nbtQEtUPpZLOOHamoonVt/5FyaxVGmwVUr8G5lMHpsJ
nR4wCs7JsSegU2JT2Xah4kJXz0hBXMzI83ptjakOuYyQNeHw73YdfSCZoRTslhlxn+IQV+eT7/oi
lqYDX/0vVe4xGS9N71TPpgU/xNGKFya9Kz6zvfLQceF6oP4Iq97tAF/LWrVa+G36UBX6X5emTQgY
z2bRZot/gdDLbk5OmlG3GRQ4XPQ+u4AuQkP9L1rylFa16V/JyCfBu8FFxP43IHqFBWSy5SUlwu5l
AHEEH2fxJAdbgnqpuqA98rDMvjg/lEba9be76ZVhXPBdJ5ivgKUAqH0WAKC+39afrfYVeKKS9qSK
Sdq7p2ink7oBrMTy8UBkSpCce2PvxLpBERsY6qsuPeZddQY9rGhTKqPmy/8Pp4lvnAcTEF+UEp9c
5QXU/dU/Z5mASgGSG7Tx96UswWAM29YC0asN8RLHEHAzm8GenCDAx8lOFntIK1RGhBjQ01jdkS/w
kG0BRa7OqrJREfqrHeqw0vA4Ie7RUjHIx5qR5uXPZP2WEL4gk8nKcbLRH7B58eJwhKruOdhbnZ/b
UktsnWwjmlymYY9BSaPXKtQqXEHAtMBajnaxoAbLLRmJpth3slnYTisSD3w7b1pVNJGSiC9rnbDX
ADd/yHjH3ufcqtC4JCWC/H1m06qVo5rvksOhfTlM5vILwXmJvcNv+gRJLVkF8ArrAwkN8pWdTQE1
x/b8rFWklR8xc39yuk0iZ5WHmTEHM9J10nVDU/2jCb+McRGDjCP6SxWm/gNvD5AryfdWLLjdAn83
i43kOW8vGnbE7IXJ6+SRbYdlgYICI4s0L6kmHLjCtmU6MOqmbi4hC1kZsUQ/a2Gy2JyML2OqAGET
8WcoEOPLVh6copJJHwjyWNRaNGfEH73ZFsVZjzY+Odbsi3VN7SJoysMZ2M5uZLtYqtSdHOsLjRPB
hEpwKmdyBKcUadcbqT2W/q/oGhGLy1f3N1xRhtdtbGz7ko3KySWvSxSSK+Om8rF9NQtUf2IyqiIF
aAsCZmguSJ+sufR9jvu4yKGuUVR69TvBotUDqz+buOUL8+0eHIYx/Mh25xzSAlkob6Cu3K0UuhuI
3fjRj2x5kwfmlUj/VAnziaOlqs1jnVWec3nyOOIztXUvEpNSu/rFez9RJQkLO8KMiQmwd5hZysbp
21FPgzn1XGDnyho1MwWAeza645nMS6BJW24h2Smq0B44urgWR+Ixty5dKfrvc+PCuAEDkcJtQ1WP
cTqRlq77pMJFsEnmJM91FoqpD+89bwB6Azg5Y0xiyJM9XT77y1PVNyyG8kqFfPFqxuGZYtSbNmaH
Yo8+9ZGofr4hS2BrpzmIjHc1KRC1aQUUCbn4OsaaI0pHnh/y5kNfzJIu6/a6zCusEpPOpuN0SWt3
PFwp3Rz83xlsvJGeAT+Os+o2J/w+HME2a1hIeasn9OoOffGDuNqo644cKHHJfRZjuBFj8zrfrcC8
wKmnMolFsdsRMxcRapOIg1H4ehuzidma/yXrdzTejx3YVbPcaQXVypk0N2p0pdoAS8ob+n4B65Q8
kl+DNX6J71R6sKyLf8MfNff8gbCUKGwWzahXJNbdP4BmGVySG+KXQqCr+hU4VNwgJG11j+4Hskqq
Niu4BrfH0LJ3+mE83E0zyp/DT0rE4s/PHoOcO8CCVA27dXPyaFi8SBHD+uMjafoRIPfjuLZBsKpE
k17vt4XJCta70ntu/7R4W35BO/Ge6+AOjEPs8xMU6m1xcmv2AjsOv03OdGYfSpTkE+T7EngWlNhJ
y5BcDz7tGVL/O5HpnGQ5EPDJZBhfIJ3lrfQa4RctS8gLFzL+2VX0Z7V5tRax477njePQc47bVxCo
uD8rNdMwFxjnYn+C5s1r6B1hJtaXQ8qGYi24lRSwPDLMqptJW6F+WT9bY2tknjTtoVOqtRIF5I1g
3yEYiNcc6mfbK+aWCNcaQ2/ZbvQta8lj7K5YC/fQ04HuIt6h8UwZJcRGppY1kDfnPFZngq4XxRdE
2ZXwcASMfZ4j/btAoXqFJZz0PUxAT1SuL/DIHstahbWb8NHr0ewBHi0aD1gLaZ/3OoCjqzGA6Vv1
q/ifvPmP7ZRDMuMPJs1ez3v79T8HC5RRQzIfoOhsAMqTNkN+LfwKWfPs1Tw7Rx8W1M9376Kjln87
i7Gss7ajUZtUSV3uBmogB6FfZgel6eSHs/a/uA7CPPsvdC6KhGrEoXFfQimpzK9TaXCxRUtS9WOd
Cuz+orH9uy7gIwazafhinOEVHCOh2tYH/aP+tmbT2HYA8lBaxSvTWfQKwDR6ErV6+sNXeYY+Gz+L
SHQMdwyyMt56yqV9lGxgGeAMb1SHNM8hnXQuyJ2FSEk+73MjW2w1ao0I2mIw9UYrcSgrg4jGUWnX
0eaUv7UWN0CpCSay0KjM2n0vb0MANdP9rNNEfVjwD5zNZXK4epCeCuWBIsRmsR5coIDvb9R3uaj8
RNONVpTVifkIRSKbFN+i1biQZxNnR62COXekis3WQT8KvxnKPmsL8bVXw3pbfjZkOFGP904vGiod
k2j3DJdPZD3WT2VQPuaZhXCSxFIEX76PCmOyU6Kmk45+JcWfEgS9Z67MOFfiz0E5QWuJocvdrMce
vtKv+GUbc+hgmLSf/VX8CyHQh5z0oOdKpeGdbhJOmC3eIlMhsWZ3X+mYnYl8gbzE47oxMkI9l4/t
YrtrL33V2P3WdtAwXApWIOxoslQzKPOaffaqGrDzlC8ec+5MRd+dsKks2da2sc+6IE6vBAZ6aw29
2yhZNsKc0aGWa4PQaRSYGXoHtksXbkVfOSufwtRQQgEoVZ51L1FDVZZ+/qX4ayANhZVLR/a1Fxyl
WqdYhlUfUd1YY6cgSX1UU9Dlv0dsVN7/Tr97DJEPAt2m4QPzhY4wJfLspsgiIKFItLW4qMEUHNk9
i/ZL6NLrrAmD0pTBj2hE6IO/32OS42ejKUwyIaPmPVH7KkNkL3jRR+0uRSfscS5DmjZWMX2cAuEY
XAVwAzGvRSxYX84pUsdBxoN5idbwqCPNCtCZYnJUlyvrn3MwBdyzzf9P8CjSEpUJxu8tjNByTiP8
LvqDQ4QQvWl8PN7QaAqBz4fEszEJNVEqpqskRl0UtL8Jk89dut4Zah/v4+5XGrGoBmfzs64OjDPy
sfhQqABg3B1YnrpuV4SCM8cxU8OFy4eBfhu3HU4QyyLKnBZ5hal3X9DoEy4yqzNC+Oagf25ruHby
aDi67UqLISuXErf2KW13mE9GXkoDaDiNQQfw5GAAC3qDx8gnRz8EP+DwLSNRSFqRw42WpNUQKtiB
JafrSOWn312RoHiiDgCdSCv3ROkMeOIr2xLpCIk/WE+9LTs5jFaS3pMtj/qSHglAVgMTReH4g5JB
NjoP4JbMKCsuRgFjNBEno2G7taTs9rPMx7Es2veHGfGRGtLwgzpGhti162milo9Eh+oTqHAsRsBy
s4PIoIgEIWA/oWc00iaNM9i2ji41wAYgugWPVmXpQDMpJWTq5eHMd/Ukk5t80wgTukG4zod6uGSh
ZxeLKrRmMYRMYom4ou/RDsitziJIDQFTbE4jHK7Spxc73C5zmPAh/KmAK4gapDJgFmrys33BFqMm
4/IyIPZGCpadx/LYoRNcQE3Ii8FgyYhaAAZ70sQ4IQhDavkUEOvD6w6kOy0e/ASpIfAYBulGJaVU
/HIGUsQmm1vgD3kncK0tzl4ufbbNhLcw2+buUYhMa/GGbIOBjy8BHVNlc22q0fEwr6Dhm1awv1u0
75wJB9vrH/sG9Z6t3V4ht1ZD10Tv8tbrEqx8F4mWPcJV9yxDoZvUUDbJZn33fw71lELIu0JqP3Ij
UeWQtRC4cNPqIbdj/ZuICBI/rdukafIK+omruZcoNyx782zSGCEqaKkOpAPVZgwG2Y5KXrj9184h
BD/sf/e2T6/eW1JmqV/njLbHnQg7u7w14k27iDfI1kdzbBQ1fBUVWz7Tljlco0cUK9vSCByFlvNk
q8EYSbUOrxzxSgPyQ3rBPDDKfyY2m0fzno0NDySy3LPNyLpwEetFftU3O0qy10NdOizQeWN6dqU3
lQwX/UrcPyJ6FavT1V6PeEA1uH2Vmvb6TD1Wt7cvlPZa3RKpI6OUlcQDaFnEKeQMajWr3xoBebuO
1YpD3dM/1KhbZOn+X0ho7+M6L5nFGKxdOchdSyoZ7gq9rghosZ0jlNZgNvc8l5GpbWa2blkdewE4
3nT9uohCCwf1AUfEAkkqWr73zCrAxH0wPAMwqx9h8302QX3Osc9/ZFWlU0HnZR5zO/JB40cROFZy
BIBS4+kKM+UOjULJ/UKxzzYOtWLy6QOozA/AGGCFrgltgCEy5IqNkD5L3q3Eh6GTvpx+FkprPWTc
qcw9sMaXEcgfzLhOZTlTGWcC7SfBfpHeAVW98UAiBTaqVjfcDBhgAn9vrInmnHk8NyKALokyv8R6
UXINNML+4noUTg7ZwQCpXB1Gyk+msBvX+VSK4BFZzWb9MTuasTJ7aP1OeQxl5I7sTqhRKDf33EWl
/+8jJIUGbf7J7CUhomTfDDmPYKkIJkvpLy/GlxeLbTnd6xY3FhdQxh9UweIf4rrF9O0amRU0hT78
2NQvvTtZ5V+Xlod+byYyfBvP6NGHH6V0lxN7IEnkbEkjFycfhsAVr0GoMcBH/C2TFDyH+ISnPP0Z
cbP6chntVN9pqz6hz82JhItIlZ6BNIWiYN5QjOq33IHsNwWRJ+J6JgbzgK6ddre+lcKbhb5YTfZ8
WfjzgRI6Nz4vAFn9SskguF+3gAQN7avbrLzV+DnuKLGBnLzrkCwnRRwyTyCq7MyAtfsIonUKdrC/
67Vw4z7CCAtpM9JTKqKsgzp3nn2zdPsmIn3vjQ1N9vvunGZJHv/nLfcH3Y9n8M9qCx2j0+c5xI1D
WEAKpCFhCoUuVYpM0sp+13123IT/kE84OaBdnWKZS5PGenfdT7pkH7odstcvfileXWRHaAKyEDJx
jEef+iEwXy753gLlFifg1rP5O+54zKRE7gJuyxvNw+d6BCc88MtMnv2s0Ixe7PY56zvr3HhJfT67
nefoiBpFzDWFd6fKw237w43dUZ2xn55zrzG75QqZ8YSz9ixoNeImNr3izSF7XHXL6m+ylhxOm/rb
9ZMMLX+v9U2iAr3y6nSDgsBT6xW4ZZoQI3ZOlVJbUx6PHdWAKBIt98d8WlsUoxQ/r30sPNqCjKiZ
Np7mXzdVO5y9ZqBfZDXN2lzMhEQdils4/Zh0p3egSJBEkuNlq2xFL6x+9Wh4Q7GZ6fYAUOB2THXe
pyQqzI++6RY/DzMNs0GMho2Qp7lYtoFcF3kwKe6Oc80KbAezvTdQcPrjXKh+k2ACBNVXuXEXSBXP
gEC9sqP+1ouGPtOjkAG4rPzEOxRGL4GLMkw6WXpCcMZn1HAWnObaArQykTbAkpuy/TDPkQbaO3X7
o5JRp+6Is4BTxukWD3ZOQU6DzVyzq/gylf3VNVQap5vw1RNmWzpXgqeYwR3wFd+HjGpYF0ZYICme
MUXumSNs+QEkRlTp6B5J5xq+bZWoicvAk015XG0mNTkWP2gECp3x5GHr4dWusAoFtz83/10A6Ivf
Pp/UheX5r/cG3nfBWgiV3AGK1Xpix9vkOF1bH+3t4YGYwkr0r2mw0TIj14CDWVzb3pRwqpKnJy0O
e2I/kBj5tZr5pSDLg0ZgqQiNiGMZE58WGCYSsdrBSJG8BcMpy+PFP6tY5zDl4abxvQYrnOPW4zAa
HdcWz1cck8luRtsOKLMTuwBW+2EYx8pd0Ct2YnWMoOxrRtuIweaFtBGkMGErwkBTIoY1XF4B71hC
jmMcDvLCFexnCWq8NWWlmK/WTg+h9GQ0PMToNunJ9UEkujxW2x6XZciWdCPSuMITVbZuqJqGI1rO
z104S1Dz7tzg+m0bSSwal9S9p/fw/ws5R/M0GJmBHYuBGJ5isPr233zXFojdvwFlYgDOnw4SACec
LFT6dPzjeAdOkukPSOLnv3DGcQYkqleq5BGAQ4z2ET+6gwhnutrkR8JgTC7hpv05vOpf1zTrppFT
WAyIxN9tc7u9YzgrubZLhpVY+wGX3Nt55Zosad85bhhy8I32iH2eAqscJyX/8nU8BaLOuyW7mymz
Ifb2WWUjADG1ZpUcW2o34f4/oH7WKSdue6ShGoyPRANMWUmpjawaJETNhalu/IDoTIWAHbQpN5ef
4/I4ei+njBoAzQPkEjtUtEbHfemjOMg6Ah244U4v3xWuR8hGeDAM506gxrGTZahB4vUKcPOs74xj
+omqHNdXYQ+wjl8rjuQH2Oeq/FYPcxmNCHH6eZroGiq+OGzfP70GPD10pEi3DGndjaX16C/IkBp9
fpD1hGvH0dIyB7/HZDLF8YFOKRuEOcBLSUOy5IIUVOgqOSXN/PTuxeB1Y8LB1aqhNLIhc2Uja+dE
ZQDxVVAYxpxrO8cf04mx8HGOMWe28d43zLhoF1004JxbJhYomi299wepXEQ1TFMphhRyrBlgtzYl
YJWUUR38aX33H7aKpGFAvYYsiu8GTmCgYeXNl6CGgRFGJWlSLjNnUxRdmJ7GUY+opjjk4ssfwndj
Fd8J+WC8zovf11e/JAEMYystNKqtpkKrwaOlYp5nAjPNeWu/pKxUXRt84DMwxfAaEYRq/FR8J7o4
mva2QmODbjEwc5AVphZsIqIxxtoy+x9ZM4L7z54qpD9902SNkJ68ZtdBmEKpLVg0w9BWBOHRclgN
SyEZzvearibq+yAUxVEi6nJvaDUjM5s1l2TTVaVcCRkmpW5YAXKH9/ICsOyRWHYytqHnUCXwIC93
QNwJrgzt3YndzRrJzMTrzEe4J0PhpiziKhaFssTP0sxx9hIBH2IMAhEYmMMnNWGc4RT+9TGLJDQr
Lc4Lg2OQbQvjZmiC44tP9Yphvyr8w4iok+CIbmXek0oNNKgy/EzgjR6E4gCeKqhjG3Z1mFNmbqyt
gGr5UHNPFRJYeWj5XNCcqu2X28K6Tmnh58Rb3Sz3pK6mO1NGHiK8bFW6UQG7i/8j6L4AxH0N1Vgh
NsGZvhnIiwovjUILpvvz80XefkjJePzl9Z5iSv7vJYMYBQq2UcjIPeTsF4V2sK/oRFovylkdtTWh
f0A/gMZQpHwRSFlM0QbNDZk1Iy3iLdbT5Hm5YV9Ouv8NzdwFi7epDSA9dqgV8xHL3TjSqKOBhnc5
vE54qgYL8WGG9h1jZPsglQDKhsBYrUiYQs1pXOMXW8Q8rqVI8dajTbW49vE71IWX9V6KNCeOTYDd
d/M4fmE2CLiMXSgNk/3vhzAaR1HOZzX66SbntI/dD3+ej26rTJqGRF9+ahe2VenxPtTG99dLYv2p
JPiI5NN7ymh6grzmr/8ZA2wftkX8hIpwtGcy/gaWnB5gODSWabo6C0y7h/co/U69qxyFv9Tty+zI
20TefuStjlTPLpMgFoSpeZx6i4PtDYa+bSMQ/Che5dn2ewdHa3gEZv4rARbLqvEJ6QmTJ1WqJpB1
+LLyfZS0xvCHzy1KfwL3WLhQGFspPmY7GzbAO6EI5+RIZ+ySieeRy6igVHvWO+fFAmTXYuUHHaDn
ZjYGdhdOiOaRuWKbu1gr6GkMvpTSvJHbg+akpvfqxEX88/iv2zaKPaM9VHavbyIZKXr8oMv/ak7C
blQgB9xp2fZUBn902Z8hpS6PjufYxdzBpcOFrUH7oMBKmLZhDB4S2VGVG6DWrNZZExZTbGiTCdLV
AnbBLnQcfKpTXISXsu2qL9+Jw8KczJvrFlpjwZYVtwk1xNgaHxjojM+nNtFQSpI+CSjIZRwGATri
DCuxuldag/sbMGoxANaXlEN0pNCOjQJZlXvdK/mphL2sJL0G0YT0zxhJDIw/TYgb/Fw+r/yBTW5q
ojDTxQn++OC/n4rMyltCOq8+oh2zMXAPaIaBC9e6KG+6SePIqjTpjWxKTLTR0+PwdqBJGm0zfXW2
oe/10654KN+M7/F8LZriBkj5xWe0SZ122P7TyWmPiD6Z6RfNBK6wdoQ6nZUkwjzcrTzeFKozsdn8
y6ZKHPCpuvPS6mZYEa/e+4BDkWTTk4qskouJ3V6goQ+0Cn5KW9CYMX0nZe4G6uAdiylPUNg+mnoJ
OLCSLZw/ouskVqVKRtJVqKKaMk7+i9CsuGU7xos5ahvIWQs8kJkQPFcIIuT+RM82EOWRHmFS+fac
ZOilYpprIZ8f1bNFXbkozGtCcmdOykEXQa8xKxI1Czda9O1y4tdk7yXVdJGadO5kmuIUiEWUql9o
bpIVLkx3dNTLbQLRy9dR2USUFbgSreKOkfg5n0G+5xt/UyC32nUiv4FAMC61sb3aW8jliwgFKLjm
ht7HaROCNMgYRq1tJ7FEShTzgWlNY1FHFeW9Kq7+Qf443rFeXn+hRlvZTELNYavUpC84WlrAXv5G
SV1/W5Ft9wjZmYntBV3TKmKMOYCxmiPKtp33Z6BSzLQY4yR6d39bc7apf8lg3cGIm/+bHijYCx3P
2wq0cxzatVBzlBYyQ0sJF7jDtaTvk8bIZuSnM8WLhk8cqLVFGUW35qLSBH2D2hJPrZAJSar1MX5n
ymALuLO2ROV6At4faB0IKCxGFgvHejgiO6mIfewC6XbQwZvlQZJYbbV2WwIrjPvoROuVAizsfZ1B
pIDQyBfPECQ/PEhsdBKCLAuGA7cPJx7bqp6ZsivPvT/80zhVFVeoLoZzcezKtyKo947kwEES2QeJ
yUaB9bqOHj7yeZfxeBlz3C7owEpTOR/0oglKDtfleEl3d0d1PyxHhx5SZoX/ivdEDNrHewWxHvNp
hi38AGfPpSTx3/tXcEPLGP9ku+R1oq+7oujgm5lYzwITSBlN4UJZ9DdVyAqtE87h9V5qlSSEQk2E
QlNGwSmYsdifCA8V9hE8LZy8mpP9M67k169nCwhN79aecRKx21BsV/OdQ52wF5BLOtil2+N49c1B
hbqHo30EDntJUOsFckEHNu8t/RcmxkQHIafTREf8RDHKkCHwPmQQ3qJb778WBrtPcMru2pbv6aJK
neN19w5WnBVFW0MvsTPhkroI3ggSC1FOnomVfaM+ZJfjb4xcvp8cw+EFcUh8jJdfkn99Ajfoy5dc
gP4CsSCHB1rTCGe91wHk6ZDeXQIEizJeNEeBRSDqRXvPqIF3N61Pc3GzhZeHpFdJMBxksgoL8Deo
pBAJzU/sgpGFbn08GmA2pyij6y7CqsyXWywSApxYUx7lw9gnzdyprUkVkDzgwtXyJRio3tF/9Nsf
hNiyVkiNq+3djQuMh62NSvwJRm4PPjTEL8knvmAsdMUqEq9yvMsF57GYmJNiGNPZfRvLyZ+et9F2
DOOX0ftgKKb/nulrw6uDTt3YLVS7coxF5Ih4WwZPLhSBaEnBvcOuexbVXOjKcSLvfN99QDb7GIJL
9l8rW3G6xLGyhctmJ8sv065VN/tKPP6h+7jJUyLIZlADMyhV//awD/wHbAhWpOeal6axBpkVXCyI
l+hJoxF8aYQf94IEMLCLnnjpyl48tOmSxy/FW/yRVeFpoX/p35gqF63MpP7By+RDRwwaCla/5LrM
Vw7mNWTYsWbZDCuzdl22c+qwDAV9dj15cChD66noTD+RLq2/oYtZrURg++eCcnUs5OiEgAZLR1vU
nys1YsRWd/mNtUmI0MjZ7nQNhaL16lVEtv4tgarCumhIf69t8xjBI6DaQMHky5Yb/oLAwiUJeYqv
GeNxCpwWORGuEeHVpqA2pWRuP8MNDsb/1rigptS5YjWmVIA+Kl88uAt2Lm9aLdsTywS5sJJDedBu
JOZMwpdceZUpxOfc52freioirnGgEVESAKa++qY9oIlZGY3ByK/bLIfGfczNQNcO+nBJ6h2vbqVs
bgh5SGinhWpJvL0oKohDGDAfEahjXaKOv4cIxz4ByGjgJdvOpId6B7CTBwjqoGA4KtpbX+VCn/3l
wHWDvOdbcdeYYauQxZ5cT+kXriMsQjWou+BxtpLrwE90HsJNA9p+ShXE9dq1WRg1lapV1Rry5Csl
xPUgCUxsya368rZ4O5vNZmayT6IC8fsaTg6mhdO/6kIoGM9sP6s4TrHf1isoxrmuX32FyaVKEV/m
SWHrUw7HLSOIHEs85MPZY1/IdTBMxFa+lokAzeMvVp8AOTA7Tz/9tiSZzQKUCcs/7d4WXMqAY+/N
X4PMpt1M+mlu6egtDKC6eGIb7IjhNamHVu5THMlnu5z4jT6K46ZG4cAGBA7duetGeu7npSRx4Ktn
7IAsNObtYoR5cG4gm3jIBh+ZzI062H0ocEwn3phd5xDko37TpCBM0HSb5RJeODtQ0Bpz0H/9PTEI
hVFvZELc6ftVj5Jl5Rp93krKLSIFWhB5SSUkeXM2B2yQki6dMvQHUP9gLYasMVIHgOQaa7GIUo7j
vkdfTNeqs0l+wKt0ozcB35d+c4k/fry/VzyVuZ71frk64Pfo+BPJbe81URVCIwg23R7ljQ9DAJi0
ytYzPbUGzHtN29vLDHmdrosvENf0AA37DECeNKYCKlzoBjAAyPm4PwT1QmeEEGUmDf2FwYW2+/ej
eGXK+AMJUpixed17ZgMh7Stm496SsQBw8R4ZbnmserymV9ZyA/m/UFmIoWT80O/d54p9ja2ankXo
twDADqhyhpePAOWlSnZLEAL1IT0s+OSn3XX+AhAjyq+pgdY2+Nd1n4IjdCp8pL9WjLEhAH/k1Ht9
jcnTl5hMv1JFeXBQi2+w9l+/BqjMtXdKyFCAMZCuSzKXrPXmGWVMQ9qy6IzhV33pQn8di6d6esAx
COtIitKgQbP/enUkphXU/2xLTivNjnLKJA80B1RbWxEbR3vTWcYQ1xfIRL5ff7NtGsALzmnxImPQ
vB4TuBPInRbRdrHy5Ikyx4+tjJnEqfLuueZT5yrrOu+LoLF/e7ylBkO/cczVohRqOoItwzQbpXSP
X/lHW6TV01Ly9pBmDcafiqzTwJm4EynWbl1F24Jjbpu8Qefj3ErLa+CbN7DbWlxROgw22WUZnuz3
EOGCwvh5Fl2IjzsyfPke0RReAHXOneEE5C8+R3lXKx80BPyXWLZn5+uT8iwvcsNo47+lRbt2U+hl
MePFmx2NGCc6CPJqKUldc6RBe7JXIt8c2G4gwred5iP3vGX0KjWj6IbJXCUVAsNpd+GhbJa+D9sx
LZ0DdwOvW3slWzAlhlMH4pnl9WfhRD1JdluTHlHkTQXGCy7P3MJ4uxo2wSc6Lop6XTNLKfuhGDs8
/0/vRI5qG4Pdx6dYyrH5P8TT+iGNpNUtTsea2bjGjusDchdaazNCSAs0M/lvg6f10wZrpN8RcIhe
r9LOvFPpH0XzMkrkdkFG6g4WTRRTHJIWvwniobDTNbzoE8x8MfxAVypfSMlLGCCba1CkpaKDTHp1
a+gMvtZt1TBlajQjrMHrgOCTjrLBX1PgwdbWPqYJeUm2lfcCwTGNes6tQJs4FM8sunpQNVix7TiP
RnrF+HuZksyLse5HbvEBTwXMSflWN0MzgZPmc1a9abB6iQuNRVmx4vpfA4Ju+CVS/yc+s/DQmM5s
/WOxTeEDUyDiQp7BazpXgfw6Aiv/GSUzCvcubK6G/Mdka9C7PkGzIlKlbzbjpqvZrxlwDY98Itvo
n4JKkLfk+jcx7LBR01ihgDDgwSfLerwJYBPy1ChMkfoTWow8q88GFlRf1jZ72Rg6nlNqmU2FF4o9
TethV38GVg9e3fCZjEchSk5pTkJns+SOWRBmxm8EM6/KtmTuL+JOVUq+qAt8+T7SSjiZlA4W49yk
V8/guleNSm4uiZDt/vos9fk+iDtcIcr6v5c3hzfFkm2MZabwDoEwQa15bVGy2LuFJPemJxDv44fC
Zx1i0vsHnzkvZK25ydGc2QfGDg2Ptxins6nubsRFRt19CQ9IOqwWJ1pbriDFfqEU2JtjnBk1vQkg
mbc5vc8K28nbQb35qS1HqxFGNMCpuNNaqWNouLjbNr7Icgcv4GcFJNM1uONAzgKvBZTm+vOZvIfF
+jcELLVYO8fxnt43L/9IWG6+AiT69meNqufcq9iyAj2WbblHyLX720R3DrAxzbC+pMwXOseVN/hN
4A+kyuyWXniYT7Zl/0XiPCvqBkMHobA1LoM4pti20N/N/2qcm98ok5cvfpmv6IU8DAaPI+KRth+W
xYFPp3orhunEm6i6yw5ox0YA3dP3/R3obCIkWDeGM2P+iaXdN15CBGyjlcwJtDIO3hUXCt8zrUo6
0LBqe5/a00Y0SGp1Zt4BxowK33uzhnFFSItwjycN9VnNQWAAQRYEZblcIXhGTcrtOJzvpVvQRDJJ
ZgXzbiQMiptjBwcFsC85QV125dCWdqL2zJFAgWTa4ZAYn6Wldztt+nU0D2PE+2q9xJxrlrZ5rIck
80HP4MbKzlqAIJMYQAtULrnVqMwUmoGE1Nglumriv7btdFIrnDfCxl2TaigCd1nd489pcUFA6PHC
82FJ954BPGzWP+f1mDSdAYOaoR2Wb9jgn9Ax1wulbyTqa+8R8VxabDTdGpuT/kPu6nnCbHYpxBhX
37h2udA91Ri2p2Ebm6cfsi8ETPGKTFa02J3e8zuQqiI8gGcjDwZzsp5ayk9z/SfgYVcsOtvDJFaE
JfW7f7k9FZHk6u/LLpqApdCRaA3ImCOjEglqPAIou7uF7CLb8ByrD+gH3Ac/YwhGAR2TcXTw/RLT
DesRiN5WTmSSZ1lxVViL4tJNfGR91djjL5PKzC5qs7GvUG+02fgRQZEG3vl6Ef4qmKA5rHq+ICOo
Yhi0pBpPQgquz+far6tBa2SJsa5WzMfXks4VzcMeMIg/sKbjwOrkDd5X+wm5bFXRTW2WCtz9xInU
7rSjeayJTVurcZChNPuA9+7AMEyEho5nzx8NHZW4LbD0alpgCN7DYDTxPN3C6GvIDD0jgexSWm1T
czASfqF326Jawxv9hI+lqhzeWHZWeGwx6r0q3psUpNlYAHi90Oij3wrQ+v7semkZiDakR8UWk9SG
4KhTzyqm9j08+t6kbML7+hqkUVcEWHsRyQipQhLceR1i/j4u08zmDG/qS/7tWcdtdLKy5oN6GXG2
KFvlTrrYLGchGqB1a1hOMgYS8HdrI8SfWndLoO5Uht3KY/E/GVfpXDqPeYsCd0QCj6Ycyk1vYu1+
DmP5S6yU+ItB5+h+bO0YTQXphO/EeJOT5vIhJDTJf0E7fJeWzMoQTqHFX93iSC2xVLBqEQUXu2TU
i6ZVmZvEFvnFUjtc0r/gvzBZAaYoF731iVE/Bfn8/s7CyNcI/HNPjbrjf9FMoaP8mu+NmWdDu3+R
c2jvy6PguPkW5Ej/Dw9yY0V76V5HErZTQDkgUsbgMi5k89biFvBiZrd4GhFsPzupTksladf5jfnH
yjIgluhvUEd+yJyGWHBsUkB0Y49inpONARJx+0ZycK7t5bNWE4bLmh+FmeFnM+O2U63LeKOyuvix
xUcW7Gw2IfPqdI4fIMBnl+M+6SZZkxSrZbO2r0o793p4TIFNit+DRzatSmsffAYIeLM37Tvw25vR
MpzgoyJu9QXnntu1ugDA5QBEzNsX90qlh4LR6M2oQasf2KES+mO8ov0i0yJF/xBqr8xhho+BiX6V
+fiv7uyXL/qfaLa8wfux1JUB3KAgCPQ1RNYU0zjO6p84K27QnQq0Qrs0R9CcFWwxdum4QXgwfuHe
CKy1uE8tXr8HSv8EAL9hZQBQejYQGzYIdcCCK39Qt0vRqrmLq5p7lcgq1LAg1HKjSMMVqA018EQI
Hd18fVnhVe6BKvKSc+kiGx5tNPM5DurDRu8c0x72C2tuJSF2+D+Mz1ezEQmWCmGlsWfI2KJ+oivu
F9RTJBo+5nrn1zy7PM4nwGKQYbAQRRhqEQMe/oRnIUC/A7eiCuYIc5I2zQwG7H7D1BXOOx1Rlk9a
w3kRWHQ5X2cOrURx4ig2RZe43qwy4RIWJ7K7De0JaAnEVA5ppGAYO8ztvGIFqARolQQWIe+IM8aN
YMTciI1B3rKn5g8zTAdi02L4SqreeB0dxoUe5EIEhYublHICEWzwXs8RNjZ+NR1l07ZtpTyQXiZa
3D9fWNEJKj23syNlXwZHh9CESA59GnFBvkyr5kCPUhC/b8XH5Pogea2l69W2Taq7Eq5vSMA0A1WK
25/Q8eKcEPxk1j/N0qs2KAuiyEh9yoTl64rs2GaJC+NR8I9J2AnbOEnNKtCJ7jrwng0X45TTXiPy
gD8CpXR8aUD4RCEm/tfM3tsBHz2ax59rEJg6ZD6gadnPwsFUOAuXhjck/RdpA7DPYRx5VwFN+ssR
TnZbqmKSCHppxiVk29r6TWtKDHjoWsK/eAmqHBFVxJLptxJUjP3NuYkow29giMFxkdXkBkI2e3NX
7Oim1M8/o+NfT3jF/gafUCDTwnq6Ou4axnCxHSadMWFoI6EosfLDL6qAbeVA3JKxEOfh8ru278M/
iFbjDLLGetw0xrdUpKelhIN29fMKpRN+/e9hluE4RGePzMdsQXlT3B/+Zpb0/2AdFj8chnPkxvq3
h6+yYPL1VqO1wMjYxbCbxdCt0NLqcIEm7VNcFxpTMMLWnBpjAmcdDE/KjAMo1PCVIM1r+8aVdkvw
3o3q/mrDHkyTEq3gmFe8YgQP/J+2OVmp9dQNnBOhFXgUHwMVcN3bjrTObF7zsUUcSnWzgiFbXKo7
e4i94L3/kZjFH44SrD/BfZJGetS0wBwhU+Q/jghbWr4Vl8rXbNhM2y8ofoS+Sy7c0tfKniE2yAsY
obfSEoOEjrwYLHfhdMWf6GfnIkA5LnbkBw9xrTBlEIgucDHEaRwPA5aqa9WHxY5cE1dbHOLz9tt7
gW3elAE7Lb/Dj7yDroBMD4iYPkZoL14i8L8fBJC1koGRYXhW06pQrF5jJfSdj8X+rRsY1ZsImRsw
aHku9V38PvD0dJoNaBXHZ/1MJE4T7W+CBmF/vop55N40zWoNZmX0ElT3dwQCOiFwPewXPyMJrdde
KpHVnjmsXyOHEOh2PER/Oku7kaJmlQXRqp4+Cw02zqSkGd+0nOl4yZQieLAKtNX2mnm2h1+94uuO
mp77uf7n3R7ZCZ06j/VwOad0uvlGxDtdu99Yn1ad3RNLO4ZYmC49gKTGuU3h43rhSU/0OROvHuOH
D5LxlP5yiI8lb1KaVYrvzLmsvt87fCV5ospng3q0dKL5XExnD+6djsKn6o5vOj+FHXf/YP5Iyx/w
NSktb6zAQj7dVayuVHjW1RIrBduc4+kmj121w1TeqKXKbUb29JnSZHLzpntgyrk+93piO/jD3VOn
6MlJBt0fyjPztqEB4w5JgZGgNDMlEf2nx7IkD/V3f618qgmklUJFi6t9E+9YDgTKV4lvM8U5R+i1
g5IQR5C6kVgromhINgVBwT18NNJya2v69t9p1eGxe7MYOT7SvIi/WwMDfM2R/677qaOO0EX67e/q
9oner63cnA12HHhiQYZX3lXOKUX7njKpvo6BncJQY6gSsEVBiI2uKAGR9BektMGZI53V0vszbVww
7Z5pgHp2I6aQhcbhb9LQQFmseWWSPOR+YpOp48U5/9Q+UmSSjUoxo7/rFVEoewaQFgGDg63rf7mw
TlJOpF6sVGYhUeIDAzPJ9DMfzJEoCQT6CEb9oHhDAGjFRvXejq+3T5cmgSwFM/gfJDJzcoBahgRo
7PMmrzDCd1pfOZE0gz9GWXMLDsn7txiSmm5Is+G4G1En3IHSU7aqwWbZcZwbrgb8OW5gjhmeEENa
ZgBuQzeeAFIhIR5mxcnqDU6gqvWCIR7nkZ0NwNoMc29T4vyYn2MUXXjvsPzy/LWwMItQtU8yfIds
BcrptWsdp4CRyuDdjJZBoM5D2ljtF2R2VA24gOzoP2Tx+YQ9BWSUsfRY5AcUjyzcbi44dWrcUmvG
6G9BccWsnqyrP2Sjyh9Amwp1qJUaK8vH6cLxKuZ+HGbJETY0tv+eBZkS9kVBXQCy6XAbsR4fhFn3
z7ka6fRxtYlUieivKLQ0voLHdz08NQ3GOKZkH0Cl1mQGpCkPUyFBzf4QXP1gY5OLwJsJk4dz9Mgf
fGJ+ZmIAxGIHs7T8rWoq76GXgRr/ar+6pnPh3rg6nKrCVEfgUpbKl+6sudTC+F8TtlM5w1EwE/37
Hzz9XRuGW2iiQhmMgC6NQoYK/OhqGB0x+bquT8wsjYXXUWrbIsaEG/KeXBEKYQS/mVGsIV8dwUFi
XkoamdeZQg/umcTpfSpJhpnewe+XDoKiLp8LeXt0cMzbTF4J+r4oG01m3Ra3C5KepMJ7FGgk/2rH
upYun7rbt33QY1Z9jVZ6EIH7EiZ+8VejvUbW19eRWe4Y3sYl6vNOEiRnYMdNgDFdqnoL898yRkbR
e8PiI924cUzwt9bJxecgguN8aDMOELGUwcVa0dwtN0fkpDhHQMeZ2toliQryGZfU4Xkd7XNL9AQj
d3Mattc54HDRu2fBsQnbW+dUsiY4+sQeYYwqJP8e28dZBjoRs2KlINUrE6L5f/+xvnfiZWrmsHDN
yc9qODlbIuAYIcUXvocTSksNmumOGeDp7lAdpW1LURzf5eNB2+EhhH05NKVtwpiK1KmhPnJ0cRBB
qpNq6b51Qk2rjZk8+7wKhhCo/g7Q2BqAjf7uUKr80l62bFc6FIahfWOhH4cbCgJ7Cyqn/3ECEyXI
vx3HpZJfvTT474kUWjzIaHKVewupRbTCcQs/1aPF3XgZcNAik4CogyKfgXM9M15/4cGtdogClfzk
nA+k4FXHzYB8gi7iZjvGvwtOl3NhzuC6W6q8mYKDA9TpDkRgwvHaiRnVkKvaYPQ6zB0EQ0/5nQc4
16Zd9v58ZlKxdNYOIW6KgQfO2ZbNju2IawVV1LDLeUQsj9SaBLhn0C3OGT2ra/9cK1Qj5lCQO4zw
xij+oQinpUPOWlvqx3bBt7O8etHmC6RaphN2AcVEWXmAffYWbK/8+C//6iYfb8ChdpiXXGSt+NAB
eLQ8drOoAvgXjuu3vRApm46iArJFOWV0InEOzb9kvXEVZT+F9K3O1cw6x/qhkwXrFj5xpAfnuEL6
Z3bZfV6w0azwNDUxDrldmIoQQQMg83HQXurYyxaVhwwIN8mbYq++iPid8uU/6FyoWZx2idJIuvu1
cdUN5J9P7ar1eSDynlmEL8er8kPDEQLCLySO8cCqBI4ABmiux7Darmkvi5ApIOjD5mLSGLxF1wqo
HQbvgfD5P/xQAwegWDcvQKoWPLIFjLxkeU76cLeyWQT2gaPDwxY1bitiI3X2+GRopXqT8QCX06+O
Vb8PeWI46LqXfLREKXF6zcha9OyUiBO2240Tnbt1tp9emYgBWfAepyrPTeeXjYX+rb9SsScD+OuI
wi3YtG2KSpt+RRjJTffNSBH5PJvCamhwypsSLdp5+fms6ByBftgD0eL6IcN1zt+tO7QmqHfyYaMO
ATbmPB7I3tSdaKj2xFJOhYe5onpw9G28x0Q6OxNsV/mvf4kx05EhTJzgy1h7iy/lUM8vsytmxfja
va49Gpt3aFnyuGECQddxhbb3jOFuv+d18kkQEkOTlRZIkZ1bTEDOTtHTObipoeOxbMaHlqqJZPrA
qE6KFNpZe+A2mPGY8cH/PZ0b3654Q/0PBNAzJIcnGImA6IMl+cCNotZBhzrlBN82mGBewWqgfD9o
r+Y/TiKgERBF891Zv1Ij359ieZy+jYpCaHJBa6tf0USGT9yLC2KC7JdymvBRwxhFeukTRu/5yiwa
Q3pJxPpQKoEgKzUp7w/ikDTrV5ryb3jYKuAUvruoKUFxgPYHqHNIxx6lv9VYZuKG33yAong+RuVy
Y/F646GctxWMmI0VE8RUxei8AFNsG8LqzRzdeavx2NYzAehVWjEBh7ez1gNn4PayGUATB3h0fIk2
YcHrSfaaetISUSlqwTUDxzmOuzOjdybY0kPydoMruojBDg3A7TycdDG8OJlqlq/n5d8M4qivwRQl
A2wJdKk9enJeUmzLLspt/uxWNju5fkBXOTh4KnCz2XYkzmpyjBssu7O3W304bX6B6nmpZcr/+z/D
MkdP9OvnXAeQJA4MkE1gxvufrwh8MLKZOoYjZry2va3LFSmcCi3bRJQXv1iyTF18adbGol0NZgOh
1aSLoFUWNH1/5SR0JlPfJ7OYEB1Gm5O/oeHx7TIk9zxbdquHsvBEfErIC4dt5asm0wGQKE45wX+O
9rpvp6Y7RU48N8B99/Qu0miHhyCHVsZSu38Q9V6ALTGuEqPg5M9luUK5YYkSmvy/TeZNPsiEQ+/U
g/Q2ozMMuBPteEsOi9RCtwjj8jg9TWGJSa45jtqrHED8e76SiEIs8JWk9/aejB11WoA0Vw9eLdUn
96CayblEy3miodkMgyEZaYq9oQuqS3LOdPtXprii5fJSqvqEOHqaHBThYrLb/QeaJ/a3kFN9OJxN
dxANM3+gUALp14uivWmu+TwGmeBoy+S7NaX1Wp5/Uy0bYPpN8fjc4AzUJZhxildpCFsuiUiMv0MA
FihlZ8UeE5k4g8Py6ikiT71NvU+8oq4diE4LZWSuANoD9pFfkQck74Ba9HmLTZFhkkrCRqsR3aO4
WOP19Do1m3ayQ9pjKCfYYoYNVA32n4SEDO5PWa1axVluChFVumgOXIs7XJxrf8Nj4TWtqE4aVUr7
s++qrM6cPFOMh4CYLu4oJBqH674GemcuF4IsrC8F/2xfsgvKAoXxVZkCFKjf5oFbXtHxWQ7y/sez
3gU8g4XjFzJxdAK/bbYviwje5gJ9wEJW4nrza9cvO5WsKgQVPtODZtit86qtI8E/SM0GxQs2gZcT
pXwDqnGFgPjX3PXIS7AnzUk6w0RZyNFlwaU5nNmsO7D0KoxlY60znvHZ+HD2fI86MbssJ05Oa5Tg
MwqXMR7lhBJh0Vg7DZrsSXkMt+goDTknyqjbs1jDTzRmubt1ARWXUuwXhgy5QWe6j3H5WGP8pgey
KWXjVndXmrs9L4t45BO+7DoR6qJx810hB5MQwnqtflEBrToajesPUwAHb7i+vGehkbLjGkUWqhZT
FREFrkYaSrjRZc9/CMiWvjjIWKG6P6s20HRAjw6nxIv1SEmsFIlMnnAxhTXXpMVAVRJJZy6/3s67
CeJmuimziZbctmRnfnXlp2YETJqSo/6ztWPZNGzYGevr61GM5cfDn869lT+6G8VY6xwRSZlZpUvr
29LbuxGDi6JGizDiAcoJtFi/ykNmW9u0pmizhc1Q/GqVyoUTotwPAxm4gd3XfDKiDiib7odVLG7J
5IUe4vdMCtkWGeV5YqKfhdCO2hTxkY4SzIvKqNUwf/ayVrGLtwbS0ubVnv1woF3fcAWftpqTdx6q
EfbXPpTT0UtRSvzn5x8WingvVuOlTSaOOFurPazFgRE0afieqQUIRY9Uj1MqKy7cMOsJA+4P0XzY
31R5ZT0yADBpGrS74fOykAzQ9LuQzETkorSBFX69Q+zOM21niKeyY7mbaHY2yO3ImF3uq8RqoBjB
RXkqRAqmu61ZPKjMVuHL5jgB+b5F6O6dNf5sxYQPD16i/Jaa8DcrXmqVXyxB5anVLBRYfWD7sl48
WgAjPoMNxvBzw2FR5GtlnC5baf7+1fNuS4BV/KBBEZQasSnZ9inLzZP8LR0emCQomUiJ2n2W9Zvu
ePsC2cCBNpv9ES9ZVUv0pjDB/YuH6xcQLZfiD6X/AJwpDO5tWvbVhkF55KZPvGY33Plx0MaNE2pe
11KTuGJ07noS4aYRrZPRCGOePG4bpyIyJKYOcgg0HDGV9fuwbZn4ARY9avk7RnMyfIY9AKtDJsDV
JsERU6Sq8rZFciNYDBOpgFY/k/FePPZ2+dEoHspQQa9uBlTzU8AKYwTX2PfaDf0oh2Y66+z12RZ/
d1eXySLVxUxMqtxEDwMTi2oMbBG/SFNeHxvh5LZnyMSslBjspdeTxB5Z5uxJL2USvgjCH/KpK+Ja
xWN4iSbIEPtCesC5RDgUdFKVo3sAO+xkFtXNUI4KVXm8ld/SiszxmsF1pBvFAs4395XOfdeZrTeU
iYDj0w1oIcNij63CyF51q7S+E8sX/QuVpqE9vSlYOHCg+pdkt7NAymengtgxUDqXmL9Ko/pyh6ML
Fzd0RQwV9IqsZ6tafR+EF2PC1FrkztWuLxnJY4aZpb58VZA7DGISUChj+eJp6HVpIjS19lbyASqf
56t4R0+Awr5qhJ6xOzeir1WwO/0iLYIDo0zMv6CKjKf4IN68R5k7mNH9SBTnHx4VimostcDE43l3
mJvuUtuDpC9zJsAcjYzJYmJL+Z5rr884r8/pueonrqNqMuFbxQBWc+rpPNVvdUmghxxXZMl5bhgG
RV+JKcKmeBI65gqo7SWcK2wm/f9tIDM/4y3OIdPjZGe6gLI7YB8fjae/RTbZkF51vNw9EjxeRSaz
u4fnHwaJRxedHDelVyRCJXmDxJPIZicVCbuQZcwSeZhq+KH+Giry5vdN2wUroYQeUAqE4vXfzsJl
oid6aykQZZyT7xrOahSK4zL8WO5/le3xGA/8Or5aT66GdfWZXFwA9ni5JS3gRymxPcU1766chHZa
1JJ/9/Msu3TpYFtz+9iNbSXLbNBRkxLd2967rBTAnHyyWb4NkFuKOvrNCTsfe/HYIs2iakVPDEzI
A1XRuBKpQG8/1AtQPo6SQl6rAvM3vW9vm4eOrx84X7N4MSu4TT8JH8FBrxedG4fi9pG5aMfTAvuN
VM8JJYQ2Y3uoaQS4T4GAyxMD8Ibu10VGLrMTMuYPhEEQyfOPtJsE3IeY95ZBZ/tvRJ5AhQjwAbKk
WQbabicxRP3l+034rw/JhczKJs0sdXJ+6CWzBC6zee+J+T6LvJLV97qAn6DGxCmeWvH/4ZDoW9Jm
+M5SJzTgCR5y4fy44TCg5u3LnQhbEhRopdM+eqXdO7KhSitmOh088pXtE8fxWGoV8SlzcMGINAXN
p6RMoO7BZ2uEFWHp3eWIW8zSDjuqW3sTBgkDAJB6TNTRHYWhhQORNBo5p+5GGBmTGwYAIjRg74GJ
T0CnPnP8xcluaJ4RlccsQ7dMuLSoZDL05l8+mnJuGOPZQZkcNBtXc4uf7PEjbjy2HHgX9o743fYR
Q20ZwfqglBmHvpJHatFyqRLEGN6TN3xtZwYpEl03NBI20bbdqsjeYTr8WLqWal7cILnH9SG92Dzv
Zu1Cp9tvttJ3fHGlmmJazp2XVaan1c62L1Id+4tyQeYUzpYct0E71p7n5Vs/Z2zG0aa4Q2ixhSru
CJY9hTyHBvEezCJr6988hesdH5HL0MvGi9LygLqTbuCclaZurcSGQdYZa00QqUbF20sR/qS5E1VY
o0sQG/ZII1R7RkZk3JdTHx/VZRHGY7MZzf7zPzqMvIJQTlx949hWv9K8hs2r2/l+C0mnrMV45YEj
zSqKzKfKi9Q9naqVt4VJvBAzJCyKsu0SKzkHcTk683m//644zruVJadgv3Iv2kd6wBRYnELsHCXC
PZSS1B4SBEN3eRgUQVe33zgb0BBlc0p88aLn8o+1W0s+wzrzqGjVyR4r5ZAYJJsXL9yZLkJTcQ+P
8bcuN0VtZM4WSy23ER3TqfnrE0Rkx76EuKuUtGk3wYJ2VSKlH6m4IwCzM51cYlw3PlX6/GxaaFZw
E2wo+NZlp0lH0/x9TS9wq42AaA2AW5u0zjJZjKf1gYAh4Wx+U+kWUVyt4E2RyBSiOdhO9D9nvhNY
BsER/Q05o/+3atAaOXoQCg/gDiuuzYPrqL/wMde4Kjy/vzuVZIuyOqGVpcqp8Yj0G5XKOXDUVXzW
lf2Jjr8sMMNP8nnsm8oNNyoTJq+Ghauc1+QLl/FNhEoyfiVjf87vvLxreJ6XYPFMXtuG2C9yOxc9
aj+7+LcxSdrV2kqNFHVqUHU7idq1thtKfX81xOZElAse09H2QQAtbE7K32c/GVwxWHejvwy4v/2M
yDYjU8jovj5g8EtD+LJI/XqOpOy3ejy0AbQx54gjIaG7e8g62SRPEYyNTsPuku6BrYJbO+yph64U
u1IYPFewH80iLvC+v3NccAxbkkIr2Xsc785OluYSL7yeYsTjlfZ+lOrtGzNbm6zrbHEpOCmpNQ+F
r1M7VhDJ5BEarVuR22+weWm+sfIni+Os9RqjltxisXLxb5ag1mXWfewEgViPj0i8vID/B+1CHuzZ
4klU89EoZ8trufj27UliprrQ9HJkAmNO3NkF2paGdLsgYMnSWqqj93DsjeShujNwfE0Qe4piexKU
xkcDs+pQmcg2JrN2UyxhByGh/VC5wApanSkfCwbTx/qws+2AaRgjTz1VcxW8tCuMKR20cXRT0AgJ
wtbkXj/Iu7qCqSqzSrq1MbfJi+Gx6AjODv2mrb4kK4KxZWuHEUA+HMyYaVRyF33sf4s4tXWUn4BB
ev7AjHDNzpxAWpslLYSzpBA5Yobl15ngxUPHp2WwCu5wP5v7DzT/JAyYT1Gkywsw24+T82o+V/+/
5fRB4qGx4HZ1+4eOwT0WmKwDTegf4VrjDTa9ScsdgYA+dwDBhTiaQP8xWEGTIxGP20oSMHd7ZQlp
5IRrSY/FXhnfs3LdxDJgsfzgWKUOhPs1w/G/IrYmsZxRiNzUfpACAaahMgsJ5nRsSn6E8819LX6q
KyTth5W0C7lbyKFlMrzOK7ty8a8bDI3kpfZdX9Mb119raSzXAQFBiNTSPooM1O+ujYY1+Mwxw177
SCAjx1/qf0CB1BvqjlfHiueZf8xAQktHWACFl11f+/wQq7ZaQGNHV9cZrOs5WtjdnjWVwrETEJxV
N/L1ogiXtxoqNr9/cnudoFNyWwxo4dxFSzeEe9GNkC/Hl2Qh+cvfBXNeShfcAcgnPQ5FypwTsFJC
weHZQUJg2gAE53eK3HR1FOg10H+9pSisDwiOQMPvWMuDiscVhygDmxpw9XPkLtNVqJSf0qlRUou+
CsYrRXU9RHHhEBdaPYrE/a1jsb1FSd5NoKNsg7ulc34Uy1/OafhhtDh+Vn4flceYdjqOt5vpeLr9
WnkutTyfJjMQoXOgNgKvAQ/9/T7zuHQpyxnPYmg4Aye1hCux+gv7Z307QrQ/4O6u7w+eSgjCzKua
3aKqoqPL4xyhK7qRYUns5BdQ2MpyU6LVVzx34F2bo69qAGQFKkHuqL3Gt2cKzTYAn6Qak9ogWwVI
iSI/WeJQFjSoAsYQ/7h13+couREm8XRe2ZA/Vg7+kEzS/jbegKnvAEo6DHB8kpVG0EnidQzCAeda
T3HpBdU/Gh61P8F1YDTiDwj7cmNScpPWnHZH1HdZRaRtYzPDfOfbZNa6ztJTBMhXnu/p7Wwwsb+P
Oh1vvEJTIhbfIr933hQWtbw2UvRvSM1BtxabEvpD2BudXZ2lEsfDBD28816RHFNGpjV4zQl4I7Ha
vbUGJuLAmvyLkv9Vicb2gOVl3f9j4hwqigOGPu9WVhlbFK0VAtpR8kClJ+rq03ugt775qQH5lLiU
tSzYu/dPooRPbFxT9eWLO0cgA0dUsshLWHA+pA+uLngSEWL43CG2rlFvBRyy3wp7YRmMkDIzLrp+
GuMYGtHJHtvNMQLRvMeElQD4U7GwpAG+FgejZ8CUU2v/ASPPxhTyEy8NuRGBLb4sBFghp43fNYys
NbtknAXLV4gzVqvYfQQ+J5MejMNRUZaxSVY4LwZ1uCeXXkDPvbbyjAaI1fgXRmxzZmK9omIGr4gz
DYsWSDmQ4iUfJm0uoanJAcVfp7Yz3EssTGV9aSyMJ5L+Y3feDpLZd5rgUhwpdus7hTqJ2IQkmcOt
X7TuAnVS2mXjfSoYhzXDqxVewZ6KNFo9rEl3rOFNG3aSrMZMS7clrayJskuDknqpaDTiLa22N3DM
BI3tgo5s2llRw4XJmCNYkWwuH1ZhZeYjFw4t7jI/Bd71aB7hXKmSpEkut6Gfi5rucvqCnn8v/cgU
FF2atbKQRpWr8KWcpza3m4Hu0Dc98KMI5+tYFC1/ofM9g1nNZxkdKicPV1l84KANF8dNF0nG57Ps
xkS5i1gix4N7V65Eh75TtGy4365zh66B4utfLDhLeIOuI6WL4tK4iyxX3LKFA10rHK6Kh8CHGjLk
b6aIGwl0HmmKoVepK6hGIN59R7qR1osIwM4H8xN7LM8fI74invuaxogbeia9qdc6ODLlIL7anO03
Gannhh5XCWNVT4QTUSDWxr8+Z85SwaEBnbsKx7FJZ25k9f1250rS8/6+2VAmRMwiQ4Bv/0e0+0bb
yyfznSGL0nPhQpYMD/lkGz/bwKQNmcNzZsjpc+n5C3+1Ky/erEHukBNJQt2exC48No4VKuRbvM2G
0pGMVE+J5gGkGlxVWvxaSajEEoyPo9578FC1wTWd8m+loG3D6HeE0YPormXm7h6BmQC02xygZpbh
FUUZrct1SEAlS3eorrgQisWPRNkYLQn3uigGB2MuACIrwSFpJWIyYbPu0W68xqnZIDofzqKNDD0Y
dXvKXBRVFoxU6rEPKnKmd9MYTmlN5n0s8FXGgU1v/UrXpd28GJX1BCQvtXLeouQgQI0JI7+pNPid
mOLmbEJwXAiMuOcehIcNh31SbzPtKPo8CcxEoE2aOpluSz1QMSs7uPJFpdAL4H7D1mm6tgfNaK1Q
e/CBIqHFCHLGuQiP+kaVWabiYVF26eSIEk2KVBpFcUqwJiqbVpqi+n4TNS/sWJ4pLa8xtcSb0zYq
Xff70b87Zb+za/twfeBVAsdU2N0G+PZsqXcHKwAbT3RAZLGFGFppQwxGoBE6NRb/k2H0khLMbYDa
eZzYavhNVj4ysEAq4oD9S7mermDsxEmRhnW6L1sRuh62N0ooAtQiBrCE2BSZ3XOa3L83L2Li9tUp
f/ZEBkLjFA95pPbgha0+I7GSR0hKTLkOYecEM3oQEB3Mz+7d9ugPaexU7LKz69VmdxP0AWEq49E3
yh1BCEBA2fy66atJmsLUjxbJp64UpWkjQDJclcrS0CO9PXxECZHm1R9kPQK4h+nYFHmleoMjWrZs
CbfarhiI5+od/oGsUAJeqZnsL4I9kB7ATfebzeRXAiGDhI1dRb3rMRth88qng1e1v+IOygHzZlwp
OgSklv69p7zM/UHGLshJt6T85/1bor8t3Z9uIxbY+W07skmDFDlaS1IShcqCwJoN9Fz+4AZ9zFux
skyDXTKS+rDQQr712tn/r/2E4yLIWM3O5c1ZuQEDBdp6ytnQY5Zg48UHJxK/kvS2eJOZ00x19NO9
AbGBT/v8/7LB8SLdBySExbLpL4upoUbh5QhQMGuHLMvf4/w2PREbMnrbmLO1naqpwUM8zBQJE4NQ
8xyxPFwqCW8196gNrvEbqz6PUkngfu1+A9n39qQiakIjMpZuYSPHoV+teM7ka6NtsnJltg+b3L7g
leAZsm/vFpwnmT1thI75adZdVp6pkS4SqhBwPm5BvF1bqwkAofJj8X2mo5xkqi3RWvXhCdjOiYj7
2GnAETyHOYKFvs5voLpEqNjp9nlcu+bFCG9pKgaEtxbgp61jdrDNZahfX0UBAhE2LjHi5wGDt8ev
TBM0gQ2YQscvnP1764a3vzMJoUqB521NkrdmLeCVsiEtRfg8pIzeMNS9Xd81gFmS/0ZpaeS9hS8Y
l63aqwz6KRCCEjpggIzjT2pYAMy4+DT1TCM1cWL+q+zLsfx+bmc08Ei5Z/MvSa7QBBYn+FHtXpQg
Uotrpy/NIfQKGk+YFREDTnt2PNRZub5h/r9cZJDImcMruCBAddTOqV9mjGSo83LxqyMiychQleFx
qicn9oCIBGBUxdE5QgY2+kRjc6bQYX42f2bFi1tD6qPu/qo5qk6pVbwtSCA57zpezuVOUJMxqFQk
8QLaGVoCcnQZpf3e9lo6/LS/403IcgiCpAPhnBt5o9YrSt/R5rg29uK2XyJkNmGH6qBsArfZ1Fjr
UwyZn6NA8RTHt87jY36DeFhTzJH9NRGqeFaV5nmmcodVj4m9lMT/bMc8RsW1ftuxkqeSSOfjDORH
STSSrY3/U2w4bFPV9etHI3IO7U7XgEu/jRXLg92QsV0pKlGle86pNnn7dXd3dnLHpQHPzfUpXJa4
3aPWCUSQEOfwR/BhNlpN2wte6GMULVWRpWFzMqPhTTIhawdDqu8b7kCcAWuPVjeVa06H7kpxbqVY
TwLZUJt2it3Tp2Eun6XhBXReRG34/52YeTjm6JP8FzxhzdUvmKMW8y2Gm6LB9EPBEMBJJeJmhp7I
Eda8bOovQfGDDBYw4YO9IgQYsvewMNRRZRlGAMK3wFdNY1W/Je4TO58GKIlcgfhNOyc/MroxRREW
jTpq6zVRA15TrLuOhnVV1gER0BwZNDouAplsVBqpWx36K4ZvM/1KwwEUw5jdXvrsyRrT0vVye68s
enZOHl2W9tPkFvCPpz34hhanglHId997QT6+JmesaCMUq8SGgkeRnmsnaaQPPIwsj1Hf5/ZqSDsM
6cAYJUtEQitg8EVBvVdj/H8YpKGGaIMr5inzEVEX72iWf1c4hRsgWq68gNN6dnVem+DxizR1aBbH
WlABAgzZyuo+MV8qNxYKVr0/H3zYcitvirp74IzNcbQzcYMjqrSze5EtnfufY9EHpzCOL+0ptVu2
UPajR7/8RPbV0BdAAwkFeuFMS1l5QPbB8D5J2rofcfQiki22LLT+uLvJD9FBnHK4jCqG3eS5LICL
vig9ck6e7PSk9ez/jU9DofDcHTZEHHUz2fUgHlkb8RAn/doKs9MAzZNwhRfvweLvZvPSbWFwh44V
62gUBX0YY1dfleu1peZyhMhFGVXc8HMNIT5xS7N6kjB8uZL0NFJXVS78d9pjgLvhR8gwvkaLUQ7d
plVzR3MAeU4a7qEs4eLh/WmY+3L6wZmS7tcKDjwJEFSIageMw8hLxo2TdkI3U2WAz56EfAHrIRpd
70nCMeCR+icSFDO6Ypj6AfmrPBNZxGuYwAudaIc6cI//rhjL1KCTUNauBRUVesKOgqXDQEVJk3cP
p3GRsWN0P0xsmxbhGKb805ev5U99AJfnVRb7Niev3gzLADGtQwrBjru4zQgWl43o8CnnnoAz9qTR
R5WYBtPDLOXPReztrUa87hQ3KPjI7T7IWB0fGy5tMiuaDPqOeYZTPsytwBzO19yOiPr5mqvIpZFr
Hu4sIbqpa3Md+AxRSkMczz3Hjv/zUCKn9sJrLFObIprsHXkdl7rOjhpKKm8N7p1GYqk+SpjtyU3l
H6PLWZGBQZPbRY53VLwwfuB5MNn5Yk33kc7BY/d7HfsnbfFKhBNeNSLNFWaISqAmJRMRY6PbCenN
H4uDzMMAuAnTbV46IL+QrE/buJwEd37IIR/qOwB3uCOm92F3OUyvrN1IUUJFJ8q3xuEDLbL0MvjJ
OwjmrptN5jcB87aFU5rc4zvSOBhXohMoQpZQ1IX1bwWL77EJrJ+Jrv527/YrtKd57wJiXCjQCQld
ZWebykXE9TWIheup6Lo3SVwSpzD2rB0k6AW/Z6GX8FcgQG5pD8BvHaAB1ZFa8PVK/Vz8Exi2fg0M
K1zHfKea9wJ4zMy61d3DhgEx9Fl3NpdiU/hm6giSlY1kiPiZ5ZDoz7xqeBVE/l8ZAQn03nxSvpnR
Or2npsKrqSKh/sAxQCbCYin6/XODO76uFVWBcAIWllxng65hvCTTslkTxjpxox/OBprmv8evSaaO
8qNyO5T1pivJ1ITQYxuARXGV+WYPg5/w0Qm6XGq5bGFBz+9W5Np3YyihTy2AQC6LRMF5+yhryIL6
iGgGbwics3EDy1g1VehiFiPnq7FpjISCWiuzZlhJvUCVkWOuzpdg+pnjrH4g3yqGJSPI/e3fuebk
k0PuEideq4VpwaWte/LpUAhbi6/0O1zpd8+meBW5qZMTY1Ab5RIkuivfN6I8aZYhQjViDmI+u5kp
/oDnp3sDvNMtwcgagx5I8VEceQEJ6qUHg1UvFxRzyBUxkfCq0qc4vbhiAVDo1TOWPzIeRep0VpBX
Hd6/gLgJp6ovg7G+hLPf1MKMG5fnEwbyt9GJDO3qIilDLvCb4cQ6ZFeV3azR5Qk1wTjg4y3V9LPP
/AiSQCJbZLjNA+CYQdtwGLBD0KO80om2YAn3I2rIJPIfNyf//E8MBLKnDeQe6/NgxBmVdAXjUKnX
YgxzHV0BGiuPBI9aUBy7XrurjmXTUmuO/eZ9y5bjZGtt7uhQKtZMlvRc62Wrywusuh6hZGmTF0A6
+Rh6MxNKtfJZpUfLX56SaRAeOPlyZdulgzL4B/Cnqbg5k/MLGIHzhT3HwJwwNeBJYYsYSNnHS1y4
Rln9/7BqHcmaAawUQFYXeN5btrj/49Wnu9DNytTBZdHuci4Gfto43qZESX1OmWrdG81xTz4DWqzF
avgKKpdZb9BU28YZ01erFd0+5j+HFUQDN87KqGI43p2F0eedGados0+ZMqEF6LGmdG2SZPTrGA1J
N8Qe6U1BPnC3tH9onUuhr5zkq72gJUWVAu31L+H3BBSojJJXNUqat9UTj9gbwfMfwfG3MOuRdNhr
zx5/humeMWkR9i7IlUAEJ9+gBDD6w7Sq1vNr/9hAZe+U3iIEwONqRb6AA1QnU711iHkGyodaOifQ
G+xHRo7FpjCQUs2fUNV289naXPDqKpXtFBuhnQg5t4X2qVmRWOypOICRhHut3rBsL/fhvn1Cvcn7
/4rZPRtL62FWQ1sYz5hLirTxT5CBiILfh1MZgRV6g2Ev2ZHBCAX3VjYPlth8m1/sALJPVspZJ2Fk
Sb/A1eT3R6MqVoXJM7oTPQukjkPFyMKRVysq0nftfxrspLhzNpABt5koYOHL5/84gez8fL0K6T5e
dQwNEiJ8ZJjfApaEtM5g6Gbr8yeCR0Fi5/dTHL9qnt02T2EKAfoAnHHaGkvvhA2aHUQh8CMP0mMF
xMU9hRK7ZYROQa3HAwj8qCWPKbzM8S3TSyUY8aykyigLQqxgevX/CIlETXenrvEra/u9SeVC7t3Z
wrLnJTtA8eU1sa7zDt2NWOFtGcqgI5qgkmBFQrqG20d74JK/+RoikWZxWSD7U73FGStjYX7QSMaa
UG1aH3t0f3pbF6IwJVsgciNG7ezDN1SFsCowMrLF6AOK2DIAstR+dY3eq01VRPW2AFlnMIylRgjW
HDx9IlGVU6Kf2f66/i6FfsVxbNXTPm8waYxZUGol0H+Y7ZwFa2gpR5yGUTTyIk2qPcKRtXtbgcKp
2exsaaSOoAY361eh8h/40vNJHAZCz5ED1ljIZ4rF2If6u5Zx7w105zctR1yUDBTzAg5wd7KrJME4
7hred49AwmTg32IZNK44F72ICyZzZfVz7hzMpWgmV+1+RqNKxImw3FSKtHJyvxVFjRxMv+M76Xd1
cMR1s7Op/RYTbCX0l/NZei5t9X52FSYCY5R14LQB3Dr1tb3R/y4jjpRQOE3nebF17gO8ymm1GGKZ
wSDCM9gDjZ14ccyoddzW/3x8nbnFNlwJ00dNkCsM3ywGMXZVX2Uu0diCXOvNQLAfii6zHDZFEIOo
i1k4yPpBIu/+zqf91tOFv8LJbQSOmsvnrZYm2KwBm/xeQGSODBhHkGl3igIM31vaHcjZCMsnO+gq
Y4ey/AA0GU1lQz1P4oImmcshnGidZxdt1Bjq5JXPX3bY+xcJyJlV8PsGW3a1QTuINtDif9j7/WqT
LoapJP7C0RlyCjx7lrgwEzh8/iRMjMm90wCcr0Db8A5oktkeeIUAMhV4X6FQ/lGKjvi90zmM7zhf
QLaBJqSEVUeTdU7H9PzZ+H9q/LspgM/zIy+dOS7U5kK2HCQHVMFqmKlpmh2SOa6nsHlVdvTXAO5f
RCuBOE3DMtqFcbzEJJSC7h3PzlJ93Ce1rgO64F41tVRYHxEC4+2c9yeBEziVJ5dyH9okLmrPN5CK
dnMAfwja6/hKGqWAqLye73+/HkPnKSRlFrYpElmsG71l9qV273vuWtgpqr5L56nzNqAcTb1uPrVY
azGseYmE7qnwRIfqbqgQvGnjeVY6IppWAiMfCpk2spMfIMKFPxrV7O3lTgcajHsFHNZ296gy1Qsb
u9/0MDA4rQF/RD+R+3RZKupSta8aCOg/z4hw+m4rCsbIFnUZSJ2Hic0wd0dAruUdVvFp8k68Dp2H
mbgdelOgV3Zpfc2mv+dn9Nmfdir/I1cuKm76ntaXBJ6m5yxysU5IKs3o574lOMj2CbdOxDKGuamR
FupHcQBKuuBb9NG7bpoQI9CkjLPgYQPSh2rtPmXIAMr/wRZgyTIpz381osMxvUVE2sseOWzpjQcj
nJZMtEaJ/FFcLEIJ6q1jgXZRZHu9qQdlJyyGxgW6aN6A+PBe6odrGPVqHWlqrCfI62Z1Vc3/RUXk
4RRcxwqG9XLMBe0SU2CmZqXlX28z3ORJyytdRpO/v3FVTsMKo1nVCoFpWdzjri7O2Cex63T/3fbt
eP/mhp80scqMoH9P6qXEczcW4WI1NcIKWhNxCA7pq1wg0y6oljUXVbDkC92nbjUF0tPidD8RZ0ok
9Pdc1xkm5DROEbDwsXgn2wqiIMfg9CPcl9S4386L8498oSoS0/H0rXrKE2qLqi4Yj/T2yzzq+V7K
9k30GiFNG4u8DTg4wTOqPRZGmXA9ZFR4xle/SVW5trq1GJLDl8YZcqlgE5VLjQntMKUU2q9QNiE4
2zAklYJ/W4uhn6uw5N5Gz6+3lFcWpqjNDEDtXKP8HUYm0XqRxP5SGUdT73ZMjXZX9pbRIcjs23YV
cYCfLFeFF3bLyi2peDJf48CNxPJh7P2RssMU+VdFKbSZij7e1OR6AVUi5pHmKulXZekEHACH4X+s
z3jINNT3w87n9zFN7P31ug7WGd52uD5MNRdYYZTUaD40YXnvky03Hi2eZDPOMFAWvB+qRhumifDm
G87pkzP/sYre2GtdASH2mTIrZ36zwBqMMeMl0LRhDLf+lcosYlzfxLiw5fvr53XdKTd+nMJ2+qiw
2Lj89YFO6WQm5lsTDFkuuUgbCsxggdfM3EypkiEwbWOmkvWXj9rJ2kG+7tq9hDP6vlAxIyXyNc4m
X42u0ZITBFnqSoIBpQ/WIaP2xuMOdvS14ahaYN3pCkHcQhKKoMLtzrvav6iPxF2E0VP2/+7BOh7D
9qtIhyht/Qw0SCMoB9TBPvYeHOzeY6qa/f3Iwlxzg6kfrak7dgdGPXhay1lg9EEllYHGAjTjeARK
tMT5/oOe2ZHh1gYD4u+JRNZBu5QrlRrY/AvxVH287CBbFzYpeTlRcrTr0as7m2vCDkcsdXJff/RK
lK6XeYQxC4cL6bFCq1vZ0SAyjafLcslqLSUC4Vi8CV5IUXV7KiZIiHGlgqcg+dqaDR8TMrIQrPSD
UbgkOY15Bn6t3WMU8RvxnR2atIov8BkF8EevOAulaPOWTuhOx8Xx71XacdV9HJmwqLTt92NctnsD
t3zlGdpJj8tzAPPaCfJhJ50MsjiFdY08gdG1fTQ/Qlug0iHF0mEt877Ii/bCc0WSc6O/ophHC7pt
wRDAGpxBSYwtB0dRllHytflwyGpDaBosnu5LK17+dtgG884tfbJ7MjTa3IkAvnj5an7Tp6nOTtlV
Jrh006/UWheBXrP7DWRCW6whwynRGpPcD8pBD37/iIICbCYJmNGs7yA60/nGlMzOqHUddwomDFk6
LXFBZLxg2pIF1O3qW30OIj/zgw6dO4E3maPg/JKwVO0IESEocLqGAynjuSygFqSPSN/jrfaqFSSx
VgMSJQDDghkOO+2x7AIV15bPXvMWfKqfDDvvcj3jwxY2jKMBMrDqPdttF9Y4JjX1yeqZwbp4pllq
yOvvhqABmc2fGmYwOefoJ60qtiSAlK/ICCLOI3pVKYXXj1vAsl/QdcavutnDRek4OZrhVTaL3ps/
NLZmzapEcyCFxE04rA6dr1rIYKocfUQihA725TQ7IFAbXUBB0bqgZCVFzmd797qUcZ+OnOvDPvHJ
+MfFohqVVeWmDUDQO2YWz32zddEzXMKWRFr38RsiLe1vPmHtktNesDxydmZmNnilp5GDVN7Ydlv1
Ef55KL92WPp6pbBAyXItrvy2Jl8sNhDO48STtLQoS5MTGYrmXDu4ZBc5WAmfRUV7qsXV3omCCMVX
e1+2Iecq5MwPt9+RGcLj3WclzQawNiYJPnq+f4BweAVUd0Z6uvfKbKNiivJAnb4Ayk9JjQDWWTmn
rssqi3pWj28NXcve2xqgwWCp89kU7/J3hg3iitA4HBZ2pFu+cqmPgwFez51cOL88O2XURJ/GTdeU
vjrfMWnGprtAJ+sDppwbEGzzaOqeJI10d8PEJ0XKTfs81IhZ2Tlc/yR9h0+HGKWy8qZtH2nAFe2H
TyzLDZfUFpyqX6/lbSr+0HWwpSuO0kvZBEADrEPCFgbwa5rdtSyHyI5K/vwVrawyAM3Z1mhLTTKb
4O5pmFceGsa9VBSFbHvbeRCvzN7ffoSLHtEn+JoX+soWTJAVS0gq3cnTBSzr0GZ0FX8S7FmY8AdD
KNb2YlXAl8P7JJnt+xexBIdcrnI4ilQ5x4+fdPFZ7rh8cGOyYuIYc7fTFwZxWxpU20fHp5I/spcJ
oQg4NceytvOIjZnU0087kMK78G0pxzrqWid/YYWr3AekIQkQxscx98y/tZpfUEJsZnznL4nM27yt
jiuyaRvRK1JbCnNJlxmIDJbseb1Y03fY9QAOaT5dUtgs5+o1iBKogR/VvBtS3Jy0zORE4VThTGoY
rlk/0nU4aUh3On2FE4xvDwZqKOJFK1aozm4R9npGj97Mq3AxCVX1lPTrhbCSd7KUrKdljpiKmpVU
9d4Lt04tNi6DLvh+ctePqUgNI6cuoJH8PfEZD6vSj+BFLd8fqPIwc3D7UePdTlgYbB6xm0riRouq
3l6TwnGsvRNQ2FGakLVMoHaabfcqyftm/EKmCHWUvlEmSuADeZfs6j0pxoSuafpmbHOOX4XlL99x
fl2DVkS6twcNhI1LCQ81uVeWCnlPSgJpMaB5QNsUsSOKA7aLi6ULTzTgMFIObqzB4jvOaWYzN5Ad
dhGYMC35Hh2NvTbwMWEae+z1/RT5IVr+4/8Afcwr+gW8ocevx0zvjhtERHhp3i3uP5nPtxHWdueQ
RR3VSkRMU99NKhgvlETZn/jOi621nKbSxLYNNI/PKXmMT7C11pHvclsYzZGDcpKQQlfANI3rPc3E
ZEmMd4/HCEfs1dIsLpM6kVpYioZBJC2G+EeSdP66Rtut3dfqkbIG7uU0gFf9efKmycJwkYNNdN3u
9/XRqnInNnuA6zS5mTHE4Nbpmi/CiBLknaQkHyN01PwFF0/PHX74j4TrdMFulfzyrvJJ9qxyUizx
j3LRPmh/XCWMhr2Cf/IAuEEVhvIOYflfLN1RL+Ps26uosC00G3oPzNTpOdblnyE3VRmAyPITuLyO
hT2j8CrHQH4Q90+mLlGuwV8qnlw7aun1a9skjAYQZ9gkHqCbMS/JoWOxjsJVOiOcVLfwOLUltlYy
9mdITtO9pPoc/Hns2ASKRAD+ghjYzHi1ajB/M109WTRE1GW7pJ8HuPfUOWIuVc9YrIxRVZ53SxT9
5Uru6Me5z9kzy1M9aeRaePcu1ztqF5LlboI+39uC6CgTapYy0oVzKW2IiW9KHANt7Hli3YkDh5b6
wVGes4PD/kVJKQnEehcOJzAIsXeyNW2agzsXiWkAjHdoOA31jdrOLA8ZJR0TNy13PLUv4Wsbljh4
0wX9I0OsDKghP82cXEXGHxujoWUfIu44UJbNQhNHeBIN1GibOKURomjTSRnwwTnswrWAcdTwYBye
HCPurQ9JEIqWTokpb2W76WKn/dTN+0Ivgb1POS/+VIBYrkKsH2oV7MslBb2EYUD26SwxLztArO2G
HQHBw7YUmGMuH/fzxoLAaoERKPUdl39fQWPp3fqmjpMV56IsrKOT0hOA0UssDqgnNtdDzZNEN9KQ
qug6kJB6Cwe+hFJfoouguIVvTQHv/ZQ6JY0av37hAnjs/D2x5nHnp3b2fF48nGWmyrrBpKKvTPSk
KBfOjSgUIHvzjWrift548j+3SAntufqinJDVYHuUm2RJVFBrINjG7Lghy3WS6XeE3lZ/xB6f0167
IR0vbiH6jd/JkNBVOGvxFSRJKy3+ayEOIyIh4smL5gs4RQAqV+upKqSBpIqRs8hZVTKj/Iu2sWT0
14j65goonFGf2c/tufLRJLqrlxJl5psOfejQGJYIjeiXOtlq+ul5hRrGSjy1B7S9gVnJk0QVSqe+
PVIcfhTutB4ABI8/fX+uWXPePyepRkid7iU1W/eDcVD37sMocDM2ImvJz53HA8vJF7FUygZWq0yJ
tjx53rA6nxp12WP8m6WizwRSjL25qivpb/ts2JnwXGmudKb6EJ1g4cLo3jLzx9eQDQeQMU9ex5eF
8NAG9Ak2TO3pdm01f7LaJBqr0aV0C9gBlSfE5fwPhXLtTi5yg2snxUGGSkr692NX4VB3b5FkbPbl
s/hZx1yo3GMag7HUKLx030nXcg1QRFmd9+Jvj29A3Oz93IIWJqKIWZ+3CUWQd/Cp0Fs37/79bfz0
0wxIHcuxqDlp9HugT0PrKhRqh3i6hY9HSRv2gSHfJzeoEtR5lOcJ9nLot6Qg56qFrMUex5LVhtmG
VU8XXk50sxsFtQFjXp33WeM7ikVN7inM2UQ5OqDaSaGH0+h6sbzAIfEIie+G5cNNiyv+4LnXhGLc
VQWxM+/bhbG56xHPSnoKd7VGA2HA0AcNtqJQNoIdRf3MVioHDE6Oq1ZBNhGXETJIlwOWKUwLNazT
+YWVpNGsI300m3bIQVP0qQ3g/TevUGZGNDACtvDjQVeXkG+8jFh2QuxWjlB4i03Vlcix8coMKCfG
lCHf5/UA97MVfVc9QVDDOyjNM3YWqc7krO+Aa6FEfYdiFBTaJ/hod/fRIyNuLNsIN5lMM0Z7hxVt
CYGqHRStSBKBy0EA6BoAZo8RQSoFHfgVj0jOk5EvY7J7d8cVcG/JM6Q4qk1S44BZsjyViICRimFj
5zzsbMlNxRfqmAYgLyT2fdxFch24ALcnl68Tna2JzLLRMI/hf4Tt8cTMmHTtfcE1lv4li2PDSYLf
dxUObwXfU24CATl7LEbbuPwsIhns97QIekWOmFWHcbjZ39a25q3XeQQn9+62nA4OsNLYxrcuOv0P
rKsDSVWG4Mh6K/1UfSXaTd05kyDcpytZCPNErm3PS8r3/SfdtUu3dANFFvUwpIdRoJoP/jW0OqJs
2HbpQfGu8H5qZUguA5r12iwTkKXylK15DWzOvDF1ulwtLOgI/CEy9SYTNVOAxOzIMW3NHwhzJrhI
RzY9s4KD+8z8+3GgLsyv2tmTgxVFggnvYdhhSZr9qAAA7YMJWk7BTwvj+A4SprgTAXp6UdXW7+S0
qdFDk6esO4PspyymrceiMy+W73z9pqkGtejmcVv33OI1gtqtF5ilJnvOqznblcUrhVlgbOjFD1eb
ajnBLhLA6+U5MEhPJDqgoBop/9pJDtk5pi/eyEr5lKFA8n4Nz56r9+qmf+Qk4cZgTjjGDE7swrNJ
Vvz9RCxdstvHwWeG/OobO8wbXfokCJnSQOgvM9+41wcDcZivo22aSN3aK45xo+OuMd0UwSKxIKFO
NDYzO+h3pV8OmSej6LimIYKDVh1nffVPY9pJkJDb0fN4v5c/OLmbbYj5i2QA4FxEOZzP2UPqgoOa
a3pMghxipv8OR9n0IpBoTetEWs974td7oZc84M1wGN9kif3GSO/e96+xb4pdL6GcnIp8VPDkI0UH
gEjoq9G9OA/Rmwrs2NduToDDDCj+DNzq2IzwiULQtlu6d5fIoQdJRmfp5KDWVy9kCJJ96bfTHvj8
WdET8srRf6T5inO0q8/iuNC1nq8z5CaNAeQ//T19X5JzuKB9z84JQDl4T5FNSU45oBvtaQHVMQTM
iwMzxvNia1NKNdJJw/vIPUDmZ6UdqGxr/bWHuNwfBel3f0hAldGLFf3AZMY1lt4Wm7ja9jpt7c6g
eFVDlCfClRt4TtSk8hMtDgTtVzAsWCbrNlZNbPJWZ62IZZ//zbUvTShGekdYCXLA1BC1YMEwJD22
ykU3ikANnEUJA05ah3X5eHJXuVMYyDHVN2t4yfmtTAdhRfg7nYkSCLychEK4IhABvjGqfpIXoOg3
/zTxxu/PI1NdedMzbUFTUxqSjwwfD9UqICqGUqLTlHnvYuRyGVRPlZBGcAAfcEizBsO7nWVZQple
O7F6nngnDFQhRnl1FICM4KJp1RppMnPX4JnoVpoBBEAcleb6ElCY1P+RREwqAs+DA/qSsxo/fnQU
dDyPyymXwGGcu4NHKzb8BBb6cZzh6iRrufDBzl7IPrmoxoAfp7cxswq9+Q29a4Td/jrjS6cHUbqG
qjRKUqgcU6asjVLtOb8TLjq3LQgRJ/xG0HgEsVFCLYSZ0DWJDWhhN+a62hvnV8r2qyLnDDB+EGIf
842RelOD/W8oDzgJ9veZdDEeoqaC34cdOj1ecLPJBb6Uw/u2APPf3TfycjXYCbaTkBambU3oJRjy
007CSGVY3L87Ps79qiDx7iF60r4X9Ih/IrIl9ujm6WpzfUFvYVgknD7XZeHUGeG9irvOW1hKkPoP
2hdq8GCLhIkYpoWtv4a9gd87DXzZVg8yrvIoxJRbivdr1dIeBLRSmFrWPdWGX4HSZufhPHYeZdaU
9OtNcA0M41YBplBG/XN0wE+upRpIfUVAGagS8m8FX14vVipluR83pzQnonVmOSwBoRJY9mmv7HYq
Xa61h0zkZtO/seeDTzWqbP74smkulb0+qVuD/cYHxBG+NDupEf2YZjExJgtXbFPddllaeggcvgZa
wXxWLOQhfrpqmq3WLCPOUQyDkdMJ9GyC7v+clCwwaPirWudJZZrjKAvDYLG9GJxyeQnphWisSI/W
TQVD1+5U6SFrOjHfMd4RNUA3MamLHn58ec0+93bW4X0X+S9ZB6BlAzZcBCbK/iDKRy93MLue5jUV
lgdDrgXL9u3tLMdGP9TFm5L7psA5Rkeaj9kCGVPx/jRZz8B+rzLoMZLrNXawhoGfwudaTJqc/AqW
m2sKnRCu1bqdWmDq3KdTfo5+SQiP8fb8WvaPVBRKHTGmxOVCfFuh2dkxGneO7mUTCc1O3suUQZb3
7v6O+4YILuRqda34Tnz7qUuVMuiYRGpMkD0WENC+v+vriEnBcqbA7dbzlnadffF+VE+ZcSarC23L
YrirIe1mvF2NYQPIYL57EnrJ46DyyodK1f4gGI5zykIlDsWxSQp4TIoNPwEsK93MHUQUq9zIGV7s
3RCTvt3qaB2rCSfHwkdDBGu4JNqUgF1pCDsyyymih4LWHtqRxvW0A2y5tuB2e4qeQvY56w9VuyNr
PGssqVuOH3aGdP9oGGmDrEsbdjfuqZVU5VjLuism9nVw0cFmpbCzuk8fCYlUcsBQBIFaK8+KLnHy
9G3/DAa7nMyLoKsLYM1q+nKLbkQdrqW17ZDz9FhA/z7UMAfcH13mZD0I0SNY36heoiCSs4HXhC1Z
l70ZSxSxS+c03UzKfoN3R/WZZP+jvSmyUH+rAljnAMUuzbfHwj05yfdKOgH51ICOZqF+8QHeneDX
8g6VZ7/ZAwrxM/Xu139Az8GrXVXR7tGyXOBjhtUr6a1RsDYZFD5Uw3ASvhReV7AeTX2AfUmkiz1c
svifFJ1JVQXJqggEImFXyGT4jyzG+tgbNZD/CagKx2QK8ZgridKx2jYMxHoyuZSg4gD8Jv5YM1tO
Cw2Ihxzf1dh3PLlqpXvQRbM74J5NzTeq7929dq4ZTBFLXBou+hKMpJYingyLOxWF3byjk54J++Up
3T7a7CKV2ypNUtiGkVHmIqsQhHGU34/fnsochtt1Hvzs0AfolSy96+3MuidoFjX/NugZ3oAR5DHq
ZzwFrPXIlh0/B8yrGqHR6fTVX8fZoqwBLVPgnxMKDJANvbrZA2jnc4oToDyscNehINiK8Tx1mA7h
q1lNwdL41m7/rPkWwTRAl8B2xtBICkBvOaFw1s7NrO0LhmAerd9i+KvivFAKr83z3PIZ7s47gRkz
dQAEmB1Wjxfb68NUgh9Pom1W920uZ6a5c+Oc5LnLRvEF1oVFu1OUlSaGKvZZPTwv7r94h9KTRaEG
TBAXizx1nq1Dg7S8kAvRVm0RzapSs3VofSqC0mj8dK9dEtUHK2vs2NF70ij7UU7b3Wgh4kRNVoJD
EOwRLc0y4UTP0xuMFGLKfMWXsARpPxnSKO/tvdecz9A2lnm5+CXQnKd002DUdvUagsLFBBwK+2mO
VEWjtUfCwybmbVj5AgtFFslQdVTcr8jaQY2DS+YU83Cjy0rrhqFKJ+bnqq7VW/zLS5xhJEhAaBCV
g77gZyNIrKITDAWTy6oHQCzEzT8NIsxxeMDA+YJL1Uz9B2Bre+cqYFxaoLpMdQzEXFQ6lzmOmhb2
3ZsHdLeSiv1LHo5T2/KMG71rC4M+pmXoPiRKieOitTgYgg8Qh2OV2LMuNa3CH47QfDswxjqd/bje
fiG18dEGXGZB0symdqrAT4e2+lKL8Gmj34gw31OqE4ez0qr2dkCY0qxIWowdueIRIzHrtN+mTlVK
dl9S3ZGrg7huokBQhux2xReCpqPn5d2WCBXvkLOi6NswT43xQLztvutBNLBNdUB7tSbv7e8hSpx1
iPgJlGIBN7aW+GdQGcdH3MS7iSGphjvdmtCsNaZ5FD2VQBhG2seWpYj6clo1zp7tVnoEgZbTXoIg
2pBQsjzG85DM4HcfBtBTxLpCKbVfw56oTkb7AOWIa8o8kRjob///WmyuWA68t5/78wWmLnXbI43/
ngwsjqnqfTVBHXosuXaRnJAiZ5XbBWf/gIwVWzDe3rQe1r7DG7Kt2Ys1eVVpI06kVBZyIw1ifdrd
c9zREctqUu0P/RE+wFbed9xoiGxpdXmYcAei+38Exl9ljNKuA7cjSFmvC6pQ6Vt0JogncFAOwa1p
FCRRqFneNaewIlb/KPt1OdjjcNvwTCBB5jiyWIHZaEo9Cvmnd8deeVWShg4H41RjpqmvXWqQalA+
qGL1HNDk32Z2AiY6jgsPP1lmdKPS4mABRJQWbVcjfTiMY0r2BD5SfN0SIciMDMu83U3OpBCXArfS
D3HovvbopiuFr12+izrIEI89VEuwpPJyKgNKpBGbudzHbai425RLW+zYw8gGEj7qQa+Th3QLoP23
fm09Np45Kvi+s6Z9ZFbVlTcF5jGEBEAo6D3P3Q15p/8TlCb3Q5Rmk7qbC+ys4XxwKK5oSBjWTniK
rWZkWoOChz6yjd2HGVKFQG9paXI7sOrVPyV/rQZbEAJ1E95mpnQFeH9QNtUW2jOJvUNUg8BtV4l0
GV0Kk/dZ23Z9+Bi9hMncYEEqdj/yynoGHNfTg+HnEWPTbU3EiwmkymsJwGXMAt+7+nP9ChEpotnc
4Qkg8a1QAk1T3lCWcZeH1fnGL+2MbZ0JKciLnfuG2JhMDvBQ/XF2120csvJZhekCYFJCecebbFn8
Kwq27qgKCZfrW5/fJMvDhbrgEdTUzCGK/ZlWwW14Q9zaB9ZgW5C9R+d45e663R7HaAqlQikCloqK
GeMcuVFZdaxC9HpKRc12UvST4064pPrdJ58a6CTa+udFOh3HDjISXwlxoN+AxqvUOQfSt3RtgcrW
iL8TloOX5bgN7L0O+VfBaHwyTkAh+MS/Q9RDEsRNJ0cc5/ey8BqIjq1tRjTLDeNbrKvM6imfpSVE
V5CypUE4V2vo1SOh2/RqdmAHA9hDt7TXitYIZYm3/2p490di1mD3NZsnK5/sVg9ZC++aEfTBsY4Z
rpNlu8PVkA1i4zIoqXTcB2AwSjo1HOwR1Wx3wyOGKA3mKRaTViT7UmmsRF0AO8t7+8j0I6V/+5wV
1crgfB/UOthgJMXmlUqc1USq4G6H0vm3soPVt+qawLHCLinupdwzw0Vi8Smjp/a7QNfTODEwlUEr
kOfOJ5UBIN0R971LnknoCjD37GVc9OLKUODlx4Ou3Aa8yRFjKCNxGfgtROND+XaBGxBNqR16nV4W
pfINNMv8FVl4jzSeKG0e7DaXFZ9MmFwizCfMYD7pSEYRgI5AcQ+6TRXWzuEgBh6qZMAV7kUhQzve
6cjFT5V6eHPeoFVHAHVLHPKg035sbgX9xqVhi0RPqY2fKX/ZrvCXGY8h3WW5qShgdisZsshh+j9i
IDhJg4pX1VOJre+e8sbGDrZ8e5Vi34K5PNT8B9lqiEWlgJLJEUqPHt1MMNRLBtywX7D0I1fg6DI8
1Fxfp9KaN3cz/0dIXIfijRPqcLVwxBjs0cN0m7fxTFxamsVTaUR3QY+rT0O+kNsyZ5z/nJPOm3vw
D5ryuSBrS9ov4SvMt4HvpovZgdyV8REo+B9B6F71bElkBuQlFW3ODo2a9iIvXTpNL1EqMfyP69kI
l+9xp690wKMABGw0BrY4GowjCWclVFkGBb0pAMsbbp1wwBTSvAiUEKXLoAA04PKN3WfQowlbcHQz
5aWMIGYonk5SH6brWqmssbDJaFzqnZ0LJq1U0k9mFMpYKlgpFdX4Ryh55EGjGmfLTDu1YVQkzFRz
zhOKenMLlXgJyxKeimyLH0X51tMT8PsRXNhBswAMyIP++kmN6xeBZIvdHVGDQzfJIKOyitMe2gTQ
YD93xoHfUXZvd13UVLau1bYtz2vt3k5xMvdehXjDxZIZf8Wt7tiHjHurK63SqZHCdgKdRkjEq9zG
aM5mTIoZgHBnh/lYtCe66sUYnJehtscJcPwSHSjBVFZ3RFiJOf9cGyV1C2U4Qn3WlmvGNAx6IbiW
rvJKoRCZ5DH00ctUB4AMPa0iYhkRVHqKE6GrJe9f4LEVHkqdlES0uGxE81OZcHWvy/L4CTQVnaML
X6yfPHYu6PVZPaPfbw8AqtnzjdmrCXySJB7qD/NJFvSg6BW6lkmWnapKJJA0ZFVsyi3lStmbo7S2
wzlmPNfKtena5MydTMwGuftpkL+FDx8H8IML5aVUWMT2+G9lUYYTjYxACNy1QmXDSx5mjc+geJoo
MRCX7Jif5JG+aAk63vt4U8B6Vyrxw+EJr1oa2lGKz65mzC2ipu2ExxDG2VPAfFoxWtK4zoR4xLyA
6xAQ2SDBuAKcGJc0vOJNB8YjrwuP3jSjJ6mxXtuBBbSSBd3cAIdal6J1GfIGKtBgHzPINn8yCl0f
VE47hWgm81RXRaVdYx+iY7SJ2GZgK1VDD1WZzWvMaI+XEAs//JCD05D3ge54uyHh6oMluGGMGMMu
zq7ktLhxLKrfpdZz4fpP5EGs3HPi+1RC6C0vvEHpLaFNYJskMxqr5SbT7sMnH6PeR/f+1flvxS3m
EbdzKj5a3J6PCOPxjVXzQAu+fSjlXR6h+9SgUi+Xex4nKUivuxWvK8j+c9pOtqV4my4IfP1dA6gM
AZApgxILubaf2gLZmm4L6Q0VhnrAbMNu1emtuqYc3HekJwJ3KvxszRxmTuKT25ogz1DjmNfmZQR6
HIdZNzJ34UiZnw2wTT+So69mH3VIfIrquhNiPwUQAcuMOhS5ZNrXKG4KMkv92awuhvHSZ1oeMyse
yNxZwVTY2hYaPW6prXa8MyFQvgkmHGUpbCF4/NAnsrb4C7jigbdVJXj/JCSNBLLsUQf4SD+1mdvB
H98YqbgA2JlI7G3r2jRlK+hFStDof4ns1KjddC129469HkChariH6xJNQ6azi1385qiaBed/Mc5l
AL9itkci3qAkNFWW503TOgjrXTVPy35MXLjJK/NLvdao+1VBZ3Q8RO9vjZQk33GhAcdsyb6DR4qF
gAs+RcYWjhyqpHA5IXc/yLY5H7nPY9eva8nwebwuAniqRT0GdhKM8zVPshGLdUS+CCJRAPmte/YT
afThrB1XmUk86viEGMLxGxpNOoV5pYHqgG3bVuW4JuzyELz6s1vgwmrnAeff+ASm6fcLmWjkgJTz
dtuG1dWBzyhAiSOklduQdX1L6RzIn8P89snlK8W7M7XSl38sRJ42GsXPIquc2Ap3KIM/j5vXxqlv
sTOxCiMDrEoSTUXRWbL1DwohFy35F/9kCLcYUI/0ljjWe2DIVpBzRJkArMHvXt7rKz5X1raQuqy6
3IzEESYeyNfjtF62C4QSKFyiMsiuRayk4VmNmo5WU00H9bwS7VgtyY+ep+4rpdFZ+9/UD9j4jo0k
ucjUVQgUij6PuW9pS900RIFJyCPN0wclDiN8OfGbS3sm19xRIRhWm2zPI7EI8mJaMQIhCiEKYxnT
T+AmkfWpkzGjoPosOozn0lnzdd4eLAylP/dydkRh65FXCF+JKGJ+SanJS4RYQlXoi6mA+t152Ouj
iiYJEe46sihtdWW8KYicMV5fEOJ6gDShGojai2TZie/UrfQelA7n8OOTS/ehLe6dGGw/PR0Tc0ET
9nrMKA6ox5MeOP3CmF5Y34/ZRSYU2aKrRHN7RBBHP5Z/257g3h65Kev7HjDfaJi84E/JM5BRCaua
olQ1Wa5E7i0dlByNVKBuYnXcYRMhLo1R9vm91dC9CWmhP0SLc/H0/e4r7Zz6dCsVjKxy4KU5fNGy
upI5ne9XdfyLtptBDzyzlgphOPEmqQDnFfaTZB0/6XsPqypNQGU4H1COiJZPFGn+BkprNV1AcK/g
Ne3cFK+xB9qN9Z41Ou9p3DC+SVyH04pdWuVe+ct7tPj8ge5R27hd14ZpbXlr9gouLAmpqS5B3K14
woa1bWS4OT6kGoJzI4D6ZccERAbwN46rkdJmUXM8oi9gqRyuG3ZZCBZpRszuC/JfU+ta9VDuMlI5
k5e9ymOgAvy349jxr8+2WXB/GzRaSMSGTBWRwNt/r6tpVWcfdH6KLovmBTnwzAfEc7IUBTo15eqQ
8vgB3xclsHQ4+qHvjIC9NHHWvkXPuXQcBn3QUJM4h9Sw+yKP1mydlIgAqi6KnqpiQd6wAcs0AC5e
tAUCvlVtTdnNZ+aCrmoBdGFROA7mXKFExl1VOJSgcZoIBKXvooSWsu0bmZ93+Ip4SroqYzmwwdl4
9RD0/ROIs9eduB92wUZ5ZyJbNEr3yEL1T+e1faR3x6PvvBwuYz8sTsMM516qYfPVKuHHSAlELYx2
l5QGE9DAm/UlpYmLFRfPTJdfyLe5qgBQlsh8M0QvLlVgnGEWcUYy2jU2VNksFMlZxTMpH6drkjxF
uEDu5NeiVSv0p4QEQfigP9tk5cy6SxdWrUu/ywl9JzYBkBc5RyWD2sLHJPP3hBvrSR5X9ZHGC+5l
Ge1CKzhm3O5NvPJqw2uMbytpEyAtCecOcFqSZy4v17dJar0ppUSdIEoGlfJnI3ShoAuaz5zoVQYg
TSaYAs/gSn/mhPxPQVKg9fzua1tiSgmmK/VjyVHJEG9WrsQEKp7/qZlWp3ibdLBb1Svc64bBKGGk
+IzR26uVr/h30/YZIfM8whlshyuB0+3SkBu48ufnZBSPWDCECzgybvz3/MeOQQM/oyWFWUl877YI
yPDV3cIij7XRZZJ88xniljp/Op8d1bWcsSmLH8l4Sxz9fQVpRqbOo/hO2jRcsJEl42OgcJD2K1+r
6DsbmaYf1XzNx8kXKVEWBZ7SQ5rHmw7V0wMjmyXUUL3hgPS+vgHGfr0ER/HMNAeXbc9xek95Zyy1
13g+dr4gea75F73XH+o3ETTKmxpGZYGrCdPAxWf1dmPgLSMEs6tokqUB4APjWdNxztIiLAwzd324
CVRUMOgb7xnVs6RorZhWN+DOCwYAJv1UTutxVW63++QERp6HmMDxccaKS+Rf9wLAY5cGcRuONAfU
gGPsdJ+60XpB7EocVshElydJZ5Llw+YrfKRQ0i1OE89P9TP3m4Dv6De+I4ud+auq/O+8meTLmxM4
2oNIns9r6psG4p81X06bDBxb9iIX16nN2EVHw5ONVZQCiG0W60tVwRF4sY9ciKA5hitKJv15Kavo
dZ0ftGrt3Ob5YUPvkGexNP4PSmdeoSjPfAZfShEY6kve1QkDM7kIZ6sX5NMKHboFX15/DwBuMXZk
PSjhaApJAnJK+/sXGjVePrVBEB3Va4R54htUkBkC5OKcyheVV3300oBgjbQaM5qu3SBN77qdkGCd
thN256r62Y1g1GMQ7xbg2iyHxtImQz3ixn5R9GuKyO8J0IlGSItXjo7e8dWF1+7gDROj/Dv4Vw1N
iwTgDz7qhVamM9zW99KDIOE+y2HZ4oEGqw8KOxfcgfm/HXMUGu3jfWT7weXuYqb3kLiFdrxZyj9Q
wnwvXKG5HhDoTI4yBpJHeiSub9Sg+VyecBGFgfmZ0jiQOggK3G3iarTbGF9dH+d4ap1D9s5JS+9a
Rpwbz3KqxlpeIZVoCWKtMfSXr4S+T3UBQe06Hia+htTFBrBHZ4ne/5Ue5mex/8vHyM1ey0EeDm+b
TEAuc7CyKTt52tfNj7tWF6y0/VmA5iAHBMHCyK+3yzuVzKBnXFepn+Pt/1Wkec8NwYf+229u6+4/
GvDw9hky63pO1dmcpSqmRFmL6qtq6NUyUd8ZR1kZgX5efR2d8PmMOEtU8pyDp+fAix36J1EvtIB+
SVw5SaKPYb2NnlL/9ywt/0a9SrM6hY9Sx9Azk2AmlmGqKYg6sQsULZzbzLeZn9dwrNjjF4IqOr/W
XbiMBqPjgcioNYExreV64Hw1V09sXFI22nmboEINtFnkpPaNAFAwcS2aPUnskGVJW079Xr5WRcbU
ix9t6MAu4el9rdKfIDMGlzjcesy0FyqS/vYuwdQreuVfgjWP4rOJ9FVHK1CIwAhr9RqJ6kZBfgTN
j9MuMb9/A5T/KqNjrTbpBAX1xfY6EW4b6Nu0nZ1HjRrXs99E5GqhHgUbN+FSl0h1xgwOkNVIe1ye
RAHDX0VnkqR8H0QNLv40jx/jTmVwPLIOqgj2JQKwY4GAKK2+GIaMYOFJWRHrKjPMr+2Vf0G/U3lR
lLdMtmlyKOJ0GudBcAaT8tVokGUEZGquwfZLmvSrEH47NjXXxzTE++qZvuhhPZ7FmJrO2XvtURFO
M+q1niPy62Rnp/E7Fb2pj2+2yYC5pE/NLReNHHwjKjIEvcXT0n3nBBVglrPSctMlQiU+D1b+nGUo
bXj3KhUv4iy4u7SptLcCQTPHXKVcALBjWOPhfl+uQeML0OtNxxwX+f/GuHdA1YbVn1ww48hc9wTD
AZGP8/61RJFBI/AloraE17Ld9KDdel9U9wVTwvVJro9pTuxYESSnga2R35z9qLZga37cquD8ghgp
aymE7n96JeWa+3Er82BG2k0tsNzMVIR3SRzR6kGUyEyoQSQhavRExt64fmE0KFfPfdXgLvfAvr5e
xHFqEqOKEOkLruupXGAw6gwwDvt9QWlhh2xXjI2hL7UkS0Q4/JsXxYsMx8A7cFdF4uGrjW4JeVJU
hBy9LtuhPTu81s2ZBUrUOgVSonAwV1XbISpKOdP95oftYPBl0wQPchE0TD+F98jele7/lqPK8KlM
KqyzHYMxLMhAUOc+L3xTC63wQeE5hqHeLI0BWwzoyhyCy2fJxoib0w5z4DzDRLyAf/mi/okPTSDQ
Ye9/rzYDwtk0zQcQ+Ggy1V5g7U+6GyTfy68IRebJB9YvJCZMTpqKjzDx1SPytQqbpk1Ti/hzC6iE
fkx0gcEKIx0rFFfzENnG80m6W/rOCS78oP0vKj1YeTX2nSWFNCpIBrsomEG5/v8po9bykDmt8g8/
SqLQr2T/KEWp6bEMILzieGEeHnU6WzP6e1dbaBoNG7Sv4a/u+tV65ZN6fkbFepLqPHGrPgHRyjoI
kfzrqVkjxKjyUUwizL6Pd8Vu3yx1b9NPyrVYFpFYqeL+Sk3gfTlfHSFp5DBA4uW33zVBODITls0N
oTJuT+boor6rutLDyAoeQKTAPRQVzh3oXiCNp2rQlJ5r6Nn6te+5qn/6ojFxqCVuNqTg/aNneVZH
3bxp0UeesfjM9J3dymEcqWIN7f4iuvaz8Fa0Te8+DAaB0alfWr+cXAYBwCDtpnetvlU3tY9+vR7H
nC6q1ONbh2IhaylU9xuwdyeCRlCuYs23i7vNIVQIf2sgpu9Wvvt4cKD/JRVWVNFx53FzGRWP5Yyt
WGDIDAPElyUeCLiLSp7Evzy4NXvtn5v/31+vBaorCLIek6uVFZpZC4wFxuYdFkDz1phUUHIX8CNT
+hgnoQR+89HGucewHZ9J+gw9k16ym3oo1s5JHB172qA63JyqS3EQEc6ziHYzfm7Lec2Vtnsp72HX
HHQmQitHN3yOb4FTTEYXjJjyfzA4m+VsTeIblbSYlE6+aIUsuMRTwp1QO+AIB+JNHd+r20tIWlp2
WCZQhUjovJzO5PYdPVDQ7f8rBUlD/7Ard1tHxHqIrtZ8OMZor0BuCmdEd8ZUzFsC/bR0wuO/wCHD
IDaYJ/B1ap7XKhpITXNG8+Jon/1ybERX9K4IqsaWYfC72PbUhUGN+ypp4W0U/nuO7/tyxGEA81jg
4KQZXzFTLQCSpGPx8q/4fiV4HNSJy8gNlQklej1jj9fJ/EEOWifraectve37wZrpYm6d81+GOZO/
0L47zANyds5DC834IzODmHKSOYuRsXcJXrzRU1ryAyG94lcqTNfcxg1RLtYuqQmzk+GRJiMijbMW
MtKl3iL5EBQJ0FoEjZt+l+tTwB8YroeDeRDAI/krCF74eAoeFs8Fh6yjfqpa4yJm1/6jLwZ1Aig+
AstEP95ID6aPieX+55ELe7oWNab4anr2WG6zGm/Pt3fFZ4dmGyI17Kj2UjKaRQfi92haeKqBfoa5
Gy1UDAM+qjWAV24cKmNQzncl6lFkuqyyrVFfN+v2Gs3/9vSP6GskmyeuHDwJiYyw2wMLSwstRcs5
qDWVA7sODCPsNdNJtr+p97G4setDjCCWBNAMj+ouJgeopjRrvBny7M8RRJFpt04Tu+wLJ3i1E3mD
8aI9QmwhV0WGgPlDgQADT6UD4kCvgnOQDK3nAIBMCF+HkkhfG3R0uTTxAQD0RdI+ce4oZJj/rbf+
GO3G0/AV3zSYrZyKi0eT6AKvn+0w2eRFHpLBQ0ZMeLYHveuEuUECi4C1bnKCw2dYFe5FX4F4UdEd
XWr/Wyzd5WlRxKE84h8PrUNXL5VICUOrfpnW6/y+zQhNFgsatuEiqu9EHG0OcRNx46QzQCq2J7GT
qHGM0WyAgUxkZeflCY/wGY4OVYKXCVaqu6De0w+WcfqdXG+d/T5XjvXMOqXLve3Pj6D2UMggvoae
ELNXdsI3YjqITqaQZSGdk4Zh8TMRg62bNpMKTf5WZbHusydaeB9bLdjlKhYOptMA0Jyi/eC53m9D
aBVaB3ODVbu71yOJ5E2BwUl6Tu3nSV43CNk67NUKzhdvoCWEukLAniRPnLA9BNapS2qnefSX5jKZ
/iwOUvKnmDN7oaXlhhiurRP1BTjHV/38OrH95esnePrNf+iyiAZ7fGD/b/viXv2BQVI2bWeJ4lAi
0w/IqsSBFCl67rzqt3W/rSmB+2SURVaq6iL40zf4IpAQq/LaAt7jAtzeGFoyeeXsq0qEddjAy0M+
SkWZi/4mcc5SoeVnYCPWOs23EnohFAtqaw8yLNAqn47C5i2zDoBafEDpwnXEQGx75XArNcjG+0sC
pPk8qyTGbEnqfO7jvAdkGn9i/iHDLOETSZQrTyrzIJ4bvHO9zoktxUl3SpDkT2VpbwG27kBt+ioD
N9VksH8rQYlNC2SvOQtGO51RCRsEz5be0IzNCH2m2QB3LChXom8lzmsKQdDSpgWA8kJty/QD9lwO
LYNhBANprmz7BtGzJR7D4luDFgG0OROSUpHWNqGXHcvUU3kwzDFqawLf9+YQE53/1csigv5J+9ie
z1K3dFJydjhn2MqbUQMJbO//Fje0pWKDzVT2nIENNxp1PoqmcKePQjokp7vDbDS9UUmmtYHV9z05
lJEHDABhdWMVxwko9uQuuYmcEcBTskZPeGCjlkvKA5Zcmj6AlPFJdFYbGpVaBSO1PC+0d3oc9CZU
dIiKNHNElmhwjAXiChBVQDGT3SPRcrpBPDuq77QIbKGyKPiPsNh5t7X6Ceb3wsuv3FBf6/HRBLUZ
h3HqBYX34OMGB8OAYS1wMdH4sEwkv+Qz6FGLEFHeenomfoC7FakHLjfINVda1OYS3gS1jqGkoUZ8
70dkJr7m3PXJobp7d/IaEwbxo1aLDmdM2k3Qo2SCUXmSKWDgLQLagrS16F5aFTsRUlGD1JxnQhuS
SBWgenhh2DpJtcR94aHf4K8gW/W09hhK3zwkE/bjUhNX3go27uuVt+3Azn+kRsDfltVmFl+8/+DN
qVYMw0irQn4v/6WMTsJjDrBc95RUKomNLo/SFL3MT0w0Q3ILnCkltlYYraduU9DXu+aFz+sRNPPW
04aFlQvHywDTJZ7EAp5tpETRPFmH3mGQPOUm+R17rfo5uuiOvNV4av9QIhrZO0mB+7Eqb21OTCOZ
5+SVwmLZfOGChq1ndUoYckCKsQgb+uxxOzf+FSNNf7lmS2qv/ibeHyvZkumMKfGYS37P7GZmRQWU
lzRkcssu72YvriFLshyr0n4ezooTfORHkgcvpKV+KnIFyHWGFi4F+mqhXOpGj9OTU/rTsRG3Zap9
MRhHK3fKCjIs5TKVxMc+x0izJsYt2FvaTwl3QSeRpqfKvb917s0xHq3ELkQVIgH6p5xBWDdHSHso
E8UWy22v0RDGWrl3dpgCw+JHmVReH+r5Lm+ht9URktZaLSpaS8O93BkLTXOaPJVWGgP0LxCs0t+G
q+kt0bp2g7diO9c5Dt3JW/LIKHjbGiUlgMMcuHVngi4HbuTpcWtJ4+AmE7SfeIYSppuBigQZgHPs
/u/+0G0OxYZi3+hAeLccd0FUUadzUcq4ExMXUxz6j6uUgjJtWM//lU8lSw+ynRYyi50SxN2ebJ2u
Xr6SredSAFWNCpwQNS2UsjbxTSAzyzooCTWRc7hx0alQM206NuLn7ci1vjWsg6gDIUSE0bZR1f4o
0UU9UUst53OXGJII0JwGkSwTe88avRE6SA8R07SwX1S4aZIfZwMv/sq5kygoN6bi+A6H159Ic74A
Oyf4aSIALuBPKbwjAvLEIRd+81IZi7iJkpA6JUm9cbz7E70IWXkNdKewlBrNmreRQvMcIXtuYuEW
NuyMqeJ9gfRGZOudIAIxXo3Jp7gQ0G7NR171Imptt89+QLl6sCFoTgQ3onAHsOy94Y+vPVSbCODr
NPOL7X9Ykm414YkOqwi4uiwURZM2AiOFapyTsVBUJcfoM9kwthkSCiG57quCxRsg3Wy0DM31P54L
HZxLIdNNUxrpc+kZ0iX0IArAP3XbIc35vXSVVyBMKA+W7tHHHgnqfXTpuyXWzBgZKm0ZMth1AWeN
EngozqXkcnO69kzYNXiOPex3sCfOmpBVQ+mUq6J2laaa+hZGl73NXIqSeuKi58fv6uEWgN/VoLd2
U+f5Dzvov0oPadeBT/W6Ki8rAU/KjtoDiuUHQ3U0voXz+7Bfzn+MKbytA3ULK/FzPs9VJuOuNL3e
hkW+Vg56+m7BIjRlssQsmiuIBc/dXkfOa8StW8g7C32DioeQy3KZwgnxC/V+8G3BE9YrcsUvGnG/
sBbzKL3SHn4OCHu55fiWXVAA1sBuvnmbt9JPFKdi8j/PLXy67rZm6B22tMR/rP2CLlWGkagkFIMp
dSm5kgpThAVmX3W3meYJEGvzr/yy5RljJC4jffWNo4M3SXEDbZHWKbfuqs0nEjMh49nlabkeVGpb
7rCq1UNCp3P1aBD8KkluR1/BRPSpDCaX1+5SphhjwUWWM15jrOgGipZ4qJFa/RHYlrzOds0czcLk
sDbTTe8ph376BT8Xd0ZBN9GNDFgv2CE6/ae6ZLvA2PXzxs54W60vRLcW3pG8lugzunp7CePOnmCJ
qA+jRsY/meghsgM3RMdw9F68kcKqJmAc2+ZUOj0AdPCcyYeX2NaSCx7sYxsxjBg6TfzWPTkaezA7
Em4KrAvzkkqZSRFlZ/LbVcy1j2o+cPKvcmfvkdYKccLxWnZBzLo9gxWwypnh0/i7H64SMtSl0i2n
EM0zL75hTm55gy+xPFNG1sB5oeVn8BTkr6FwLHZvc9X73myc1IKuWU29rZZpompBkN2KiU0g2kAi
+20VzLZTVUVtil9Wywd55LzYOkO7PNb9bq01WqpdClNTpRxruVcs5J+tTagquo4R+xlqgyPov1vT
01xww3x8Va7TfoD87SBu8KPBZR/STDflhtewh1yvLo0A9ng75Y13uAd9N0jY7VLLjusjS3dkYCOO
85mgNaLR2BazXUmACqAnV8ol6SLwsut0q1zPdqs4IktXZ6XQoSGpjMy+GxqKKz5tHyhuKHkfEko8
/a93yEz9fMslAGKSQlJ4H/1+13O/4zt2iR7vqrdFWfD2f0MilbevcWz2K9nN64LsA/lgiEYv/Czu
ITMu5snsQ5H/yZypN5WgjFjIFg8u5wgjyzLwK522KqRKFC75R/ZDWSvQrs2/Vr+m9n3Tja1Rg+YS
s3csoIVI61bfoFlfkes3RgxizGqXWIGwn6xt2+7/6gFwqiak/VgXXwUBefXubG5sYzUGa0CVN5+v
kqcHwlOmZem33dBkbb3tgVndKluzan//olYWi7KVAQglm4OEltlB2hCkbEH+NCQioTPPGpfebhWZ
ZlVkXwR21JpO7MsaKAP3amy59lEZOBa9mkQ+z+M0vVSU3vgM28mrbu1qU/gz0ZkTxv6LywDYK9VA
2LUnH42k5s2EcuycwIA1EYq/mJoT84+WtrgNf47kt3DBVD7s3bcqIFXWHjWo8jQi3Q94dENY7S7n
i8MgYRoJoV9JQL84npsk53WjzPAz1Quz7aqf+iI0/kNtnvbbR80uuIDSuCRu9rNoKFcTMnnAE8OS
Tx+GBmuRDJ4wE9OdE9KlkUf9OZ0V2WJ0sWfo7lPcv4C7w9Q/ZCcW8P0s18kTjHQG+fHOc3repO6h
/W0HKXx6l7rpKGKdW/JPNqjyj7QltrrzHWj9x2j/jceoGYKY8J3Kg0q3g8Pm9JtK2//VCk4SU5Ft
fyehipZJSMLGuixOD8bmsL6MQxJKW+pwDRCZxMfC6u9YsUS/AOjORuuecYKvBhJAXWFgNdj3ceJa
hYjO3OyVtwtmon+VNr23FEGBQGwjM1OBXZDH1tWlvQqq30rkqVDOaNJrzHk92USOONO76ioqgrrQ
XGMIGVw6WZdKcJ/bVpsAEYP0HUWYcrke9LaeeCcuwEnApUo/uzqdu6EMQ9MhE3lam5wLTMPoYyVM
wLpUfCTxzjAXEQBuOPB/VW2HH5sBE/mCKTHU/jJxCWO90rfOdXwYAK8/CqVbEH+tp8ZjqfV3PZEc
em7KTSt1MhpE5fENe3XvmzMURJLQP5K4ZovvMB/DiF+7Va5ha0tDJZwQnfN8oKNfMOyso06z7WII
fpulOWAunKB1eosQHrDz3FcJib19Mwg0RBoJEBGY/RWxJmnRAT/4i3Kt9svaTtJW+XStyuins0NA
pInTSq7w0YXzcHeVCH6//+HHuAiSMb/K3tqllpyukHy4od7dkwDfS+P7dshGWWsu/HV2akyw26fq
7mbr7hx6RoRN1nM2xRM1ehwUtF60S36Pth2sddbK5xXF5aT66WxlAgJa/3hx4vs3/dlVC48+aCSY
tcqWiRhkau+hb43yWHzjHzm7na1AfHng4gGj0LzP8FFHGIugB9J1USm8NqRLIC/IqPudxwd2vsod
+Qdn3HOkZHdMhcJapdR5yAjWL3voELqD6v5Gbbs1Ygdd2O3bYkg4zxeAqAdTn7xiNgHQ1Vuwsan3
WDZ9XQgasrYSaVOlp0sIrKUJPRLALzkXzdgBVt9Uy1AO+2LGzPoUjqKUrgedHWQsraQk+VS7v6K3
4Vo+j0L0f9cb2mrw5Hi9hZb9pfS5hDhmQNejP8kkwJWOSNtVb2g+5jShrUCy7bkmgI6u497n0Cif
ndgEfhBgVjU33x3/cvhwc8e1EpOVud1bxwtmV+XtrNteH+20yStVygJrtKMp9fC6Rc64QgBgTIsP
F9HjS/+23qbb02OVmh484nsQ8UjETpXV7QdagTIwDsO51WdOEuhj1iaMKYqpvfPwAvmUDQfThmYC
5a8XZwtXcQQxuYVOMLmEI+ueggdcMZuWzWXbBn4x6iHWcs5Oc/duYDY7Cweg1W6f7KvB5aAdP7YP
YRx2SI+JzhrRpTho06khQtFhgca4Q3867X8TYSWsvXOdqbbAC+df5IpqjsMQva4p792YqAJmJAa6
1skXSZ1o7gIqEj40JWt0zuKpOAZavuLhO0vHDOHxjU/K7HhhRBXSerCp/tpQJIjHNmyksdlq9FCg
Z78/H8z/LzaAVomN20/FODK4vmP1+Zk78Mdw4tqkEQxRh8c0P1TZxw2ixG9T5u731IPcm8XMgYbi
hDnqZuiNEp0x/5BkHXoa+oViOoUcAAEnY3gHWljwMEJes6kMQxCQE0f17Au7/RqZ+XAGJrYuW/31
VcAPHUPFo2Q9JmZVbMVixYkn4KP/7lDq9aLwtLdNPgd5kZEc4S4usiA2GzxZCg84sczu04V7k3rt
2C98xD8D6YUgekcimtAhwvCdTH7iTl26TO8z8dpDoNBw10j52RlDcWpdWIwRQ+lmkfxYxuEkmdwa
sBIXVhB1QDvjqMa5Zc53FYNQ+IJI0/lvvvK5Y0DZgxXfUBUQjqYA0WPAh1vn94BAyIr4cV+A20il
QX1igeJphDozgp0dWN+I+W9+i0o5lcoRN2HNufGuI5sL1R0ZoSTrV7tcYsKPwB6IWll8E1QyvuUu
TDYaw9fq5XeX0vF6+PsqLXxBTGnFfnyklcRE60jz3Q7S4f+1G/FSPOlY5+spoSWm8/gsbodfL7fV
IgqwhAJ00WGKBm4IY9454saTD8zGr4r1jhKCLmjFemuv1N19zPHkNXVpgGADtot8m9AEYbHVACwR
x78go4xjnvHpLWyeqwd40//BvqBhXM8iT9n7BbuHy7cO16gjhdnRM+HYrm+tZUujacO9Nz8TLm8v
Oz3ITCaaL95hOTo3O2K4p0WiHbeVh8xGp+wki3wxqt1aNIlBPWk5H+iyjUcWTeCiGR/0tWol1dIw
Tp52X5APO6AEdn/U1YYthxbqqZGXghWMTOtmhDH3gCCSR5JSn4PB4DykJIiEAX1jLMdabEG9iA72
Hkjx/Wxb7ofVL9HOmu522OlLzX3kl8O+SHGmyhzWqw3izpOuQc56ClBTG153mOqPpaffpu0nckWv
E0Jy6yCu11MSOED6USqCHkAxKdJ1kzh4bByijYLkvRBZ8NA5e6jS6PZw+TFNcE7Lw19Flx/kHbdv
zYE1rs3g2e+wHNbBdYXL/Ed9x/i/UJKzu5Hu+ZKAtiKyPXtMidrQQUH2YruOtL3nHrMjWIHYLT5F
0GPnFI3FUdYTrLM6+v4aCthdeHf5qQv/y9337GB5bF2ZEcAW7Z9VkQ1x9xn0XGdkf4UHhZRcwzkC
jfQ7LwJghh2eEoSTwCeYHarIy71GjPG8NG79dO2M45imbsiaxEo7x1CgR6Ya9KjOl/KOp6pBQ54j
vnrFSs1hS4z4U6hmO8RT0AptnXkkbhg07xNmkLzDR495XDxRz9Y2AH+D4ChGHeN/Vf2CCgFzfaxN
JinzZjuPKK2z3CI+0ETW1xUiOeoa3wfUsukPUULmyFlVjcO6hH8EzMqGO6elCYosCBQ9JqjGAnaU
1eV5yVvGGBZgX+Bj1ByTik6G6vz0ebewSwfI2cdeaeSSCJfSE5pVEP4k2nwMsaX06xZJJ4WMQru1
+ETKQPuOalXsAHb9ECbye2YMkWRzShtQgjcyR/p5q0vXyLeWVjrEfnkeTPAlLuh4alp0seqIagT7
qS2A8op/3KVpEoY2pjKOF2vl5bOarVHtEighe1hTQt9kGpZhIZmEL9RW3205TCuFpdFLyFoz8Bxi
4YGQc3+OIEaYrtKCXaCq3c/trWWxmDcVVbW7fPHMMXhtVnDfzIyNLEHPEVfUikHMjFMxLoZR1cQ2
/Vo3ZCQgq+ZPHPN5VDE2A/z8ieTX1KeGmEiPtcPVm8Nn59LRULNukX8FyFC74tRL9iuP3dbk5wQo
4QttxpELSqQd5phkAei24c//JpqYls1uag+72BNBqsd7XXiJR6/XKBaOM33PwRfGRcwWplJ2xbnI
CNYTCRn4l/ZF8OFqYBt+Wf+lYuduPUXNNf1CcY+PadCLzLCR07t8I3RX5ILxcLCuCju9/lCV1Szv
LNSzzXccf461qAuHzkj+x3wVX9mkTfL0fe7y3EvAYRokYVUzRHbTUuIrL6BN6Bn1uWi2FHWGqwbV
k3rRHxmNQrZzKsGXCzbb1hzdGweaflHZudnqABJzxaYbUJop3WcRaJevKaRlay+4n980L+IzW2FW
EjOJ8SQJfqYNW5XkkEsoHbXLjmORzCwUjvyVwqVIDXyGG7clrt3yDFgdAh5emATtcXcEbZi/gugP
WzRfIGDurRHZs7+EMvIzYab4uv6DoTdO5KNbTIPKtH+9dCQ9ek6CuKbGcKelAGzqeNgqtYC+Z256
chFpb2cjC21BYrqFMNK0k5EgLK2PPRduxasR55HFBZUf9jnezaJNgTb2HSIrrM7fk8rN68IazMQf
imbF/FPOy1yvMIeOM27tkTsxcVUyj0FkA5rLl9Y5snH2IHIc8ZPPHTEmeJXvbfDtVhBInCvtQj71
YFasIv0UDnowh5L6MhWuVVbmP0vTIqK6KjdkM0OyygQuJfYfvhNMlQnQaFpF1fdP/hztyufxg1PP
L21OF7EQ9CTcq06yFH2NKBeSDMyFh5R0LllmQBeyQ1KxPWBtMCJp1OaPPzV5kVPUwSBeDSauRJla
KHA4omexleQZ0+acs0Z6VFoUcwks7eF0fU4YDZvveAOglweHbnSKmkUfKgv/hFN59PWJoNIdScQQ
wx8GiKXz9YkgEmYeGFiWu8ilnc0lCghIpKq02RdBTdGCUSDh8RrVLpa1FEYFOIJ2lhdPTgZNH1Y2
DVXQ7A/YnFNTUhQ3sr5fIPQ9oQsZ2rqfPu1s4kKiqPCPd2K23JFhGx7FWQXB8ofGOazlWDSkTz6J
8TfsguN+mTrrHTnDNNd4FcRjD25hol3p8T1ou5tL/+V0jDUxANksloqBEbPl1CUSLrw5Dn4C8ej3
V3a39RgtfnaeSF75QfdveJEj4a/gHDTQTCbuwUTAswK85hRd0jwstfPK7TmMJl1Tf0s3gvRaXuJS
/KSIoUWvLqhMrj0qG8pqFEyQti2M1YaoNYXO0kDNTk8HbmKpAJapW94OpTx2C47+NvcTZXLOnk9s
i7iW/r9x9cb6lQuwjn/zzNwi+I4LorKOOquZIyN4bDcMWi0Z+lTb2WhaUsxghExMlAdq0HhsT0Im
lw/EtaBb02KRr3YNK+m9ckjlYulLAmSZl3Z0HLfUO688///Ge0HA1iM75NmsQ0d5F8KXPVJmlrXc
3Q2Rp+bxTw1t/Whth/66yV2FDEx5QwSBTTYFc2J4dpS2wwL0QuHbxdSaeLOJQvjwJn1ze5rdSpqh
+Nw5zanXzDaijR/2Q301dHQY0ZLVoduzMkUOWhtttxpLbfN0Yv/MRqa658SNv+WwugWWl0PyY0QO
2I+/ZCPdxgn9hTWFq7iUvsyHT2bCR5ER6K6IPIS0ogef8PmY09fkGaya7uqzvXcx6mGjwpy25RoH
JtpaosQSw8LXIXJBc/6DUMVprxb3yudnvnBPYsLD0WN+xuvivI3oG5GTeZ0cjKLP6+OQ0jFzFRGB
sjBc4mhjlqvG7TY9dq+GgzHN8/Adodoi1sjrC+KjP5+yasyCIZ5yHa3f8bU6U9H2hCZPfmOk4Omd
F8bzK5bjJDd6FCgNGfmta57EGm7tesb0MImrv6GXeByVfBQUZF4/3zPKpg1Kg+eX7LPQMEP+cj14
XaqKCGaBxKLnwPmnK/C2OxYUFqYAaLfv46yAhcQDKqRXvq8SI1RgJOMzHYgMmHB6T0YLcuG4tfd1
2ugRxUbeKy2T0GPtd6YT9SyEWr/eMaATtQwkihmRkmfkmJXLSpD5I+mPonWN1Dkgy/Qyu8Y8BlzG
2T8gjve41hkANclzDjyB2PTzXFLjLUMhDxf8zAgGSV6i+4frDQBgKUanPLCD93h99/Di09wqKVOr
SJW2VkUhWmkXt07fgspPBFLjG7pruNZLni6X1ZPKcdgLC3VpzJBkUR4I7nF/wDIaeL60vEHJoSQj
JJ84o4E0Ym0QgOlR7JqzTmmPm22SmJWfkjT1mQkf11nXeX1Cf8Rs7donQpEXOPFS1TEBuJHtkFlV
GuBh8ICcqDNyUlcPQw5vt1fbwr2teyoK1sHWih/60A2aP2O1JbaIn2p+GIwp9hi2gb1D2XhUqER2
LRrtTPkSaEqpAo3ANjQWkSicZHe5E1MoC8h/RtYxhEyc3E3MWp+0XUtIlUogrFC/Gbxfw9T6AbnG
iulMBekKa2uChg3Zaq5GI4GJHrj1d0wNJqNTYXiDOYObyG/2wkAaSiSuRNUG2brFtMB0up4BGjJt
Zd28qc2lOpkWh/nFfrZhEyKZ0PyKR2HQ0p6JQV5J3o5CtCmm3YNLub5bDglqO68i2ncEAYkNNMK3
ru1SiNh5UiPJ7SFShEvpPR0Ru6Oo2eeX7ZugMik7+RZi8OLRg4YHr1zrWx3mjSChEfCxTtCIK0pK
VyWlY0hPfXCIRyg/x4defyQfD6JFVEGLsdgy0HexsuVtNrU1XgGh3ZZyNApXZymLgvLlstLRlcfI
6i7oqu6XOa7lnGjX0Kt1tGon8vpA+yhhmGJHVozWJT6K4uBnNHES+1P9EK18KOK/BFPiwO575NYY
oh5GeiYzCws25HppPy/dj2eiQxYkfnO24MYPfopF5HQY/ePpytF7OSmrTDOzDS+c0LycLohRlgmY
vGXG4dL3NWia6qS8VlKVZA7PQ0WQZa8ODOmZMaG333yIIWgRh+f7Hv9ad+D+mMuf7eO6cehbEFvI
E1ODPBfeEW22uz4JzoDefNECi4LkAmnLVaWJ9vlCnntKePcXobS15K/O6Zt6kdGTUK7IIPcy6exe
F5UCxxyHIhTywKMRrpwE4wXsQK7/OYhppESWN9tDHni94DDWx8YXQKctwAuYmOfoV99DqxjSvc4C
zuaKtOTJx9VNvHDGgMgp9RkLdaGoLr+su4gF6BCuZltJg66KLm9fiVJbrHETFT+RAMvXU+sZtdrB
vZGYZ4IzJgP5lB28kv9X2Iglivd6UL50jPw0xRKY986dNKAPJ156vpNzl4bY+4uk6FoqtD7TsTFd
E+wDd8LtTo5TlNI9W3YGwwK/fCHuPbiXxXhBJsHp4hG3Sl/h2nyl0xRMg2g2Lp6nVseFpjeqOwQX
45TRKGhFl6iA+BysNa1/3z4znLDLE5+7P+wHyazC5cs7tbGqUiM/6LQpQTB3p6ij3nMh9YK0pvFb
NMWVrhBk+zB+2OodMP0q3TcVmiBDJ6JKrQ6hXFDpa60BmDA550VnIg6sqU+FiYOg0AytraE9MB9F
SXNi3xApFQ+2OgYYQlfm4dwokKV8EHDdSBsSv+0tHxQ/DztCpQWmrkgK2OU7aXGBcN8DLyG9HTkh
tS662x8DcIO4oYTy18WeN7J680im/d16RB+D+GpAHYcBOF05EYG/vL/wWFO4rIxY21y5PoKR8jno
LJxL2OBTg+v5mfeHmr+PvdfNbsRjIEhsAJg292lo/xKxfi+yk5IsxH0zlqOtfXR26l5cG6+3xecw
x0MtmTKyPzVMdJK3TTI1lemJ4VGEdk85rIJEvBGB32KMQS/2N/HOXX3S93O2lzP2NZMqkb1IK9Rq
xuLDf42yrrFslK2I4MN6AtEP4s3bmsZVMa7SGu6oKQfmtbyieWddjBFTe1nEvjL9Z49FjVNarBXq
QQMPFcBL0f3VFwDrXTYserDnDrs89mGXVp7Mtp/Ul8cCut+fqPTpB9oezKFTb2iG4ZbHAUhd1dhr
qxFPl2pQociS+oWxejZOjeUYlDKweHcAiTvl0LTmXMnFVG3XvUGRt4XsSxe89MUJyaFs8oxS0uxz
MZe6/r6SK4c0GituxvKZ6Tqvj6NiAs12jwGpl46AGc8d3kPUyNx8iYCtqVEzBN8bvxOOjhYvl703
OE9C40lncz3oc7DlIxVcPA52Pd81uuVvI44hpjty0r0gzgcJ9MuuA6ALSRJ44TFPamY4FYWXtvmM
wczwJkVra7nnon/dJG43uQdi6PjWVwwD+nJvE/lECSjFLKaVe3RUaBnGb0B9Wt8AJgntyALsy7od
iJxr/KVjwwwh9GwgPbKP5XbWfm7cmmmUn/9hUAv5T0ln3wT3vWjuAs8AaUel5chKQMTG3jhyhk/K
3AIOIOiA3ZBWnCuXYRnjX3MZek5R1NN0LSkxHeXjt6FaEHT2fwd1g/RQjgS+aF+yUfLdPqIWyry+
Cu1xuFhoxSJC6jpCfSglX7bwAKdAHTGAHAhhuXJwyRZ+VUyTe7kTkSXstjTF0HlNPl332ELudRWK
K8CK7lviwjIZ19cKx5Lo5QnANtIrVRvM3eodL+v3s+q1K8swkJh2zbMU3M3V0ZRkZHjk1wwevzSt
XgU0/pf1Z3LJy/T95rxt2XatElsjglWsyxi2j82zOxXwDAxHGIQFGRMNgUJEC60qtInjVnJux6zL
I5yc3Cs2ky2XPqLE67MOswOdQf90H8Xk/qbGl7KTUO9k4uTjgcffvj2tmTcgMNcuof5OqwSFUM0N
h52bT73WbABJ5V6xsqabNJQRfMNxp17Bht8Dit3Z8VdailjPu3lPL57jZVRqHweiCgYMe3Y8YDTl
FR1MQIduUqQX0WJt1ZyYovz7Uxq8tUyg3yioMPR+30Pm64qEBaUnWj6UipBvwj4xl3QDi6t0mESF
DZWOI3sR4Fa2Pw4L2d4TmbPeBzuD7+jQ6axlX+rCVwWm6inBxCeWXRGPo9pXHRMD9JuoIKvkmHli
lBJwQQM2VomoAvdq0AGD+0P8IqneXsSRX3CdSBJZRLtfoETPho6w/f22DXHNTy9r0B2j55rrQ1nK
a1ICuF7Pm8TY6mtMxdZJ/bjWPXhLKm4bxl6bClZSyLzNYpbvOPI9Jbr7QfHn9Homt9kPwQ8NEtLs
0EmNZMbElbIyhMI2U+Y1bYDLKPSk4w+KNrZPntSlselpl0NV4pl1PKcmyGwr4ZGeU7AYX776GdLJ
KWITJvioJ2ruDuaWUeB+7ijh1NFjn5kLOkvaQLuYuKlQWGRm/6uRJd31b677LTFlX2bOeW87iN6e
grZCfp3UkGs/QLH3LwagYD0Hs9RWpDvpo95hB8XT0ORsvXyec/CGwjgPeRlY39FZ+nAsOQD1uozt
NuRWudxHMyEGUrWz0dN3xLRFc6EhDxnHEF8Dlkk5BIbFPZJSn2XGBmlFUpLOcxSyoQ/8ZEW2FlB/
THAlGLXtaUhQCvFmWdxl/L7l6solYYcMfyh3+yYF6ZIVONKFHpamNI1Qa2yQc6AUNKs7Ns5hW1Kf
FGe5fBp4bVpmuI6eCDvVSgDt4qnrfEnRexlTw7yyQCQJ7MCfErA6C5K5xafNm3VBHZuihsWXEaqd
h6A7MB2ltFRTsjIF/PHMBuMcOmX/2vPVkptHFdww4MKKQT8wsEoKdNdYbsWerKS5OO3Ckwmo2QWW
qzkB6VTIHWLlVRkdQgrKL7Iwaxc4gOfVa6+WXf/tdngtUVnZS0wmbHiX63lIVndiBaI8qV26mRjT
Ulpns82DSzZuTnXJAoPm1zaBqq9HyrHezdOFi7PJao6/NO2H2gcbrppMaeSxPXRY2KJNvbOIFTdD
1RDg0JvRRTRej74g0U7FWHXJ+WJ2qUtGxper+aBdzcA5pNOM21YbRk8E0Zl1wueFL5uK1fKXSpKN
s1+kYZXtERqBftr9Vhv8ZH7h0Xc/gBW2FZCZBWx7iLqPlS/g8VOHJJeaV0EsoATUQtMhRu+RFJgY
ydUr7vaeZVwjwVffzcpNJQvgPWZLAVI0RBB9IhCOH0KvPnYwFAMNnHLomxjPvtLPmH6leQZpQr7X
I6ziGo9d5IKJkMXIPjBp8uLYqCdtAMLmXuycl/v/SLbUiLZ7d7JTLRvARBS2zCiTCptzHBwHLQGL
cShXRPsk1wbC/20k9nny/ZpruqN9Xt17P2mQs+I2Xt2rzGT3eniNEIDqail4hWJO+7zAGq8fG4UP
DigvJUMSjrDDi/mr5dlhAcqE9881GSBq3FcrBxsZsgtxICMGcrlYVJJsyJLMg7XNS5LW6oG3npfh
DMK9RmZCfHxf+Pe5zZACEy/fhOoLmbu7MQ4f6CVF8s+EqgzIA23tpXRAiLNc7UizF3ZD2R2tRodn
AnzNdbaTfNfLSWBOfashGrF6Ezx68tOh586RZrh4Fa6aZ7TV3MCFVeJTnVQTDywGPdRFunOM9/89
MPIeJhoQa5Ja3uiLr5oxaI//9LuByjzzoUj2jYKpbsTJtfXuYqdJ4b6oKg02354FC5/Lp2h0F171
r3HT1kxQTYAhjjsJ8tgk5YTonrqmf5q/U2WGUaJZy163i/JTA9g1l7hvKx5rsYhyWLAY0YGXDJDZ
p/jGXIPFscgJTY3lDHZf+0xHQ6ix4O3Ox4eKQVev3ZkVQ7mVOEdaGRUpWYEjXqV+n7mE8AcC47xx
GbLwH/8pH8xGcmK82qb6LX4aDfT/vr9dJCjqkr6XtrW9/8NRD/FYeVgI+iEn4/92e2lGC5ZcvKCM
+hNbnC6BwUii3iqE2e1lKu1bwbezYklfxFcdrRXAKfUw1fIiA9tXwZjytqIo74g3upDRWm2f4KJF
W8vBd1qQQkD653T/t4OpPG9IqPFkbm4S6cN8GQCeevuPQb79z6EAqWuR83T7dDR+6BLBOnjo/JCs
uBor+ccair2L79nI0PowlgFUb2IxdryM3b2AP5Tm/USFb5ucPgcmOQa/sVwhKut2cZWAvCdbuecT
YrjPvoB/QPuWr1d18ouI8Vchdg+qX4Y3NNifRDi7LDe0sDc/gU4rPFVz1q3FEtFUcvAPwoYHVhHj
i0eiD7ZABCKRSDKrEdP/fpjPUrKuNu06Pb/a2rot6FypLmi0WuVvjqdM9ZV5HuBlVm7QQoGALmBP
2wOpt5dB83mwpu0d6C/gtiDdLWd7nlOsrIp8SaIxnjTPmNbViYlczFKjxl0tPVSjceqX8UD35JMn
ZWWwHuQM1d7pTjnrObGl3yM9Hapt2fq9uyUuw9GZ9Vrn4yD57M7pAhE/+yrksNBpprqR4LUI5bpN
FadZsPtiYmLzleFCVIN0rynjNmPKFDC4WEUt3rlsd7dKI9hZFHfJ5b5oh6UTMQR24KLYtY2XYRbf
3dfMNzvfs+yRcrJ9hPYdalChh22Gf7RZ3gWo33KpvmSZXS/j2Cp/XHlMfqmUzNg6WklaKZuf6J1Q
TWFQoA+B6AaBRXI4QWpg11K9ZchPf+fduHd6Id5Xguby85PmtiPj4HMS98zXuca+XNwSZQjmAuGk
g5p9ilpUZRCYntdkuIhwnJqMhP216TSGWdix8z3zoOmK27swuoYY0oWe4MqVCEUzg67NW9GRcCA8
2uEPsTTOhl8BLXi7BZdwH7b8aB+uHMlGuVt0MtGfifIoNzUCkgO60UdRRaFqMP7JU9dMfVNJO61G
W5ejheF3NUHUqPq9kb6rozW/FOAjhON8rWmdFALHVyidTf9v4YW1m866Pv0e2H0v6GNuBxpyBbri
nhovBnAMJF6MISUHxtDuxgRizwWviwhsMNEnxwjTONtaZ0+1XMKHzs2HLB2BqgcCnRvvdZtXEvy5
pLPn45JhleasFTiGRSexkbQ9Z/MNlfMtH/NR89TCL9uazueTuk1Aeo/qpbKGqL5dQn61yGZrbdlS
tsTWbJa7HgFtGMvAVbRsGGIxTfJuR+MJEjIIPajOm3u1L2Mc5x9bnOQdP3j9Uy+0hUOSrYfYyu/6
WcuKSKFeZagdezvFKATep8vif4ikYj7PUtnBwPGtHEflhrBXdkGdmy49Q2+6yCucTKm6GX3xdd9/
hDsvTpPwyqvKcMcGg8fYFq4K9FZHXO8JBj0RM7iq10DG1qUAJL9kL3C54HJH+l01n0x0t0fjvp/p
9pg8anI5zfGmIMxVGKSviyfQNpDl+UnWMT7MX4ACwa4gpxzNcJytXfd50y8rRK098BwyrMsRTkjK
HBj/ri8xFd6R0l1kOWo3EicrtsOT9PSJMH2i7EM657tHBRkkX/2VFZTQfK7zHfnVISD9CRVwLdqm
LIsKuWIZpu9bCXdHEeWKn9NZqyh30rFEMf1/xoxFvjQWUr8u+i2Mv8PyDANMuS3bHkUatzDYyMGn
t+Mne/Cz09ny3GqGQpKbOBBaB/WFgtzNYB5qr2KFm0DsKpNVGy65Ai5LOZxs77lj3X1pxa1TOymZ
k6EPpzVt0NVGZ8CUIT1mBiwGhCqhJgb3Zh+cSKczyxbOKcM5x6yR1fiqjfCdCBjCsJxfWaAZika7
0tsR8eWk4h1LXJtFUZBa68j5b3Aykvv6pBmSiLinPr/A1Pb7u2qcFg8KDrT7TVnSMXZgSf38jOf6
PMD7WNbxqotr5YeJxKgvu7CoYrFKxobh/uGjFL7MDKmqwHzgONLXrhpODZALCqxYwevgfq8mFE8H
jOejrLi/lloN+9x/bODFDJQ3nyX2LxDDz5j6C6pf7by9TgiUb1VBuj9JQPXTU6h7ucpl5ZhNF7rL
pukjA51skcsRFd0CzhlqvIPc32abkVhxHaciDJsnnHmFJnP+adxqxA/YuEWRdPYJ05TLRlX2bkz2
SdvzhvlUYo3It4zJuWtMAomXaOb0ObGTineUUDJNQ1WQFLrSvhHlqlY0yQKYh1fWslH97xi89wQC
/qjL4EpBLUHpnrGq6kprJ9quY7a18XrLfSCSbUjFc4FxQx86QRR40dj2MlvTvtFeUk8SkoLlXheJ
iB842oeug+FK5PZjJ58Yrz/17WdCKcD8U25L2OHNOmenXTj1S1GS8rHA07vXGJ+jO/XBZevewYnE
EhWEmOx+hDtobFs2+x5gOcpEZDgMypMlBP7k0H7DwT8Jf959q1dboMsX4hZZkApej/TfvK11X/v1
qKpWrKULLJYKRh5hkvvLSpYvkKVpJ8t1TPvpvoF606NZYNyApoew5uNZEY7VMBcb6WmHnKAwPq9W
SCYYdV8rZFiui2ytq0/f2mkF6gE030QV5kuZ+GMzsx4nLmBmXPY/1AdoCx6he+gYIXuoLbgwtdgs
ufRHUYpsK3nAie5znIFEe6aZ8D5nbrmsNYLRebqkf0UbWtIraADycAP3rLYUy2uOrmgzudCZOZva
da6vo9zSIbUpIWGa60BangxWC4lj8L8WWouy25YWf50/fqtu7aZX3hMek7JON1SNHsefQYFHvKJC
sAQ4ZcF84vEP//ci5OhfeVOdm7p4sUxp6NfbQ+HN47rL4w87qupUjpaJwWdluTjbvOoKblTqY5CX
SFdSLLhKCD1PaAZOsFY5mlkmRIG/t4VEw9usDAulhXtOCTA+GMd53qV/xZngns+EPo9E4fBpTnXf
Rwxdj2yRSTXzHglu6XKzOzE3yx3L/iroyPVG+ttA4Q6/SLgzHYAyVy+djKuWhENdpkc5Y2PSpo35
PAMsDH8YinpwHdktGoYaRJxLvfqap1u69YNnE3VTlfc8Mh1rIJ5HwTOd0mQik/PzEio86FMO1xgd
Vf1GMrYxKmELPwBDNR/XbLlpqMOWzVXz6DJSbizIa8JLdWZoB9q7G3ePgRyhpUj+/gThH/hNFsb1
dZNwmwS34Wlx8jDqj6mE99t606Od5iYxyjFftqmHb/U6UR55/ttmxqUjEOGgGmPiBSvHeihXtkLz
Y6FJanM4vTc4hfNRunskOP/4aQxq36Rh312yq4XZq6uz6llmXyXfcCSL0ao5ngQdUQoBnWDE6XoD
f4UwSX825+rOucXLaCD2IeZZorcyTSF8yLTKM9uXmPVfwOGb63o+sgcHSL6yM3BUSfdimoIIt95U
j2nD3e8ltg0GLgP1xjKtH1FQ/huKTcnclaEks0BIIkLe+r/VjHtMwmlY1ZqHipyAav6wFlAxFopG
tNYfEWHRAAw17zXhCwl5l87iXU/ffPAUxHXIgQVDEvlUZSa9yEHfS9ikNaH7B/SOeJ6LUOqUZrBV
JUrdXrHzRnkhmB6apmvWBijMcA8Tso6DrxbEPEB2xFad5SHDTVZ6zVbpYgRj3aFL5JGP6FScEgqO
to67HncGs1K1Sd4osTOuVlGBsdPWVXYU7xjrgj0w/umchCe6a2pSXdOpM+xxtZ2hpTpgHQv+eXUo
Tkdp21mJ9UWu14TGp76pPIEqf7WHaf+XMGt5BjROBgIa0yRtFD37SaLL3xWinpnkd4LWWzLEQTyh
jXF4NfNVlSMj7jjopnj7jC9C8kPJyZW+m1crU1/ZsGGhEPLGDWCi1L0CCSAaIeCUouxTft4FLpLW
qPCfrYvjEwQx/oFT6IWXyEyJAEI9/+S1pDLgHA/JclHidU8jwMUlDAKiY6amlIWd4LLm5ZqP3SIP
YQ8o8kCZylKXNP/jFZJ5yf7KYIgjhJuaDanzFqsK3GaqztANMRJq3jFmIb+a+Hxb640TbFLg/6YB
8ogdm0GMbzBeDRw07bpFNLyqmRi9MPHjACG5g6gsfCh3F6ImwlS6NdJHUGYOHzvMqxdhQVYbz4ej
X+lIzGWAY2m3mG7inbcXydHCH995S6zlKALINyO8RQ1mE6P+ygooPrWdGHojod93GsQqnqIFVbI2
YqA10FqjLI50HJgbYMiJVs5ocMKjBrWySN3vnXgBApbA8TB8Rv7qe1ybtRU/C+uH90G1O0XefOiC
gYgeIr9CLchoOF32QRzEXrjCFOCZivLGp97pBxlPXuAKRv+xz7e/bKXpZQ4t+2u65UCoY3KSmJDg
KgW8OhmBPP6j6tsr4Ger/KwOhGyk01+n3NkGebcec7QFUwoFl9DPym8o1sVQy3V9ARDkyIjWL2WE
JcXUO6CA99/CV2Br2K2EKQtbvtEELDirF2VgWVP5NUqbU0J1Hi9dmMVmZJDb3teRNJ2a1WBFbKkt
l0qwfgDRhJ1dDz7qo5xwxWZO2MyxS8ioInXingz8lCuOTw7ozHPNag1u/UfLqkwlSTUooWY9UVmC
UbUbvlzZgqE0FeQqZvsrg6Gnf6vxIDZfFnYwUrV8UQEZ4XWSY90NKUQUi+bBcOqQk+5SUpPUjVKo
xbPATJpaAFS/XNPS91SwuCS2pgutP+/Fgs04ZMWbqCmhAXlEdM5/UK+RRmJFri16S1hBSw2X22To
YrawXmWFunj1cM/apqnYnMvcIPwDX8mbqdYTu3e6DkgoFJNfr6hQFgAZhML/TlIZKr01JPGH4dhV
kPVaOOJxMmHu0WWzyHdMfcVRUBJvUPIeH8gG9/H/J5Aa2fj85kNzXfXNswLJx1+/cSp8twORS9z+
PpXFVM4y5zNCC6yQ5uijwZo1ZJOiOHkxf5LJC2zJY4agMs6SZadGomeV6IsaTYtAcxikT4E9v928
0Pp77hfdlTfPvzl4dradDWq9yR2NljWZcLGpuu9vIsWEvJw7WLoW5fUEpV3WSgGTW6flAd5zEJze
aU+uZf1nms0dezViIeghJog1GjvODEmAe5X0skfTugd0bKToJxz3AEKhT7p1LTmOfCiU1nXw8hkd
1TcS1dyTlXxFTTHpcSBADEtZtWbD5KdMQXSowU7eurSm64nKJdhh63DpjDwm6WM7+ngHXA82IdG6
ykgwqKDVEZo+cnG6WJEHbMNRjEH1dgz22trr+LR0zzxuQbzSbPwjLTc0rQggvuBQoSQQggO79kb7
7FCKXUcwjU0MLVlM3C8aL1rscB239JuBrAR2us+mOpDTsBTt/Wh0GlEzgSQp2hgJiO11ITZtTH23
TTOb/iOfREvRQE+XoCWEpmbphq07psHEXGCpgCJslpHJPn5eDH8eEY0tluXVZ0AmipLDguV/ARMh
FT/MmvNbIsMUZjtmbLad4rJYTct1ZuoSHtjTpwY25Qq6cpKzuU0amtHV9d0gjnMNkFDeBOoZJjjU
RU6ceEWPrkK3DCsI3isVYJNFMxvOY15bnPG8M50XiSs/qxULw4EnnqziujExScSkb4ujZGOll8UR
otQUIKmmMjYVnmdB2tebHTOj3/GiwSnV28tiUOwYRxeQcIRi+vRjdhKke7fDyj6sXLr8mal+piQl
dw5DhDOt/HdsiSRlU1KQnCjSR55NgvmzJJQGN0xcBdSKAcpLnAHTx1lQO56wXGp4C8/SS1Owq1rI
YMosxwtrlqRR9MuSHNbh+ZTzbJA2FVlAxoyFYJjFPzG1u0wtZvzXKMdOpB6M+1hFOYLaCNaBeSFZ
WMTLOsgE3wxexiun+n8NE/MRmKBUSU2t7L4A29BK7hMQ6RRJCqgs1hh7nrqE+uijHFZOVfukwnB/
wlFUke1aOZKPpfCsgQtdfUuWEqeXC4RtTtW38u+iDCIUb9aUAMBW9Mp6Hm9YqOBuosA7fKlQwQfi
xFXMl1B1Llm+IJupnUyR/0yOnvaMFb/6G0O7keDjKpIQsCmmVQYR80Czi4adMZm+gptfYtS6bfU5
0WxaU2/stXhhkutmj782q2hLy3CWzwhBxj5+xC0RAecCUhP8uti0U7IjuM9fVWfERou0gdBrzHdE
xtvpJAxVhjCxsgHY3gVQvvap10ImfaT207E2uoaJ6iJZJOOE7s6vR2qwmQ1i08eaEXz87JO1m8Ej
7fvvnOH8NOKbGdQ4acT/HJMnZ882bjrt/1wm9lgLBe7xoePilyGN6xmTdbKY4fYd1czfGwkmC+xu
G7ol5sBC2v8uYXIzLyyMf0IrD7ZAmMOyPnNaHmR+MUYm60VmFa4XZ08pfgtO/+uO+duCsVSQOyub
hz+RMBVvFnLUgPBTCkJ9OomQ0zU7BqDZslIoauz/wLG3998iIbpofAPiohMAIUx2130mTBddiled
VUOZiQH3LD4qfGFlatWyKAAWXa2W1DmFkBEIFbFq1NNvlO1wpi0S/yI+/FhyvtxvDwbpWU4ck/yh
bWz2a4fVoLrSV0eW0k099beO+vg7r0U0FmZJawA3KqLHOFCtxI6goeAKdNVfiKI5hV70HO79riBV
bL0NuSW3ctp9dLRvKmBgac9RAUDhmCsAZrTxEHOFGsFsILC63VptrKKPxbuNaUQLwiV2Fcvam6H8
Byqfy0G4c38hDJrbD4NhbpHpNyvWA+3VRJRgp3qQjVS9dYIG3WUp+VW/+xvSrb0pdDA17FMNA4CJ
EEwzzZTIBEEAtsbsbfJdFppAKovkyKQuzdv1vZtkhjLUa3ObHfe6gp2yTtsiC1OQPU7PzsM7UxVk
Eswc87nuEZxpn+IFk/rWcmbYamA2WI7cMgmNJzKjXRbEQidLjfrEE8QHeK9gF5p5uAQnNniMv6yr
rdmW9q805+C4prYjS/0FslXW4O+Phu7d6DdUmi8bm/3szKfidkDHd/0dRqwvwzdK0yP0kTwh/r8g
aKIJPWDyUel6cuee6kCFOEcUQaeJ8ovxcLaYpB8JIF8XZuR+hhfY5WiTpKC3xfJLOlwV/KPJdQay
tCTpKKLqNIfcW0ig4+LSCra5yZLPOFZscFLsY5/YbUoeKWMmhA1baaff2DOf5QSsD9Qg5hEFpdfk
B4zFUhPOfH9PTIe/IcsC4vzEv2SqzdxfiZbJ1nffMgVH917XWRRcz+62d5ZaNqir7aLIbrT1OKu+
6NupnEL5xPLqDO+1EuDoamagJEsPKjDW8Ec3GSOdC4eelDEC6N/CyTbp9wHDQOcJ5PZUZpBpgPyp
w8n6VFQqlGXPRTXn4p0/4I3TwcsJ2hwWsTWsqPytoeWhx1EoVZDP5tFgmHOMbW+ge11N2W7SRIpM
6XuLhggnLCtqfwmPr3URD5houa7jt3qu2btjP7jr9nlVCtcuh5f7fuqdbTk8RNLSGKP2hqomq9+P
0yQkOSeRU0UWigOZVVV6BSSM6QCvNRyHKHyjEEYZmmV4QEsVt3LTSwmNRU7WEY9ayL299L4Kmfae
NdpvTewPrq91ucnpZzvgOdCSrCNolRH5XH3cduFE3E0ZcjH9DWDQapceerggGyUYtZvx8lXNyl7x
9ljwRvDfZXSXXRHgZ/UbkQrS5/PTcOs1xfHT5a0WdFP7MXY0OcQlzcXpwXy8zrj6eu+uda3x0e7x
xCCrig53+WyJhniYUH4liVZuJXX0HyeVrGsLJmseVo6rtd5rK2nuCjO+MQ6iuOpxDyC7sl3azFSD
GrrTAKDfRJnUscCHvZLHBa2IGUHTS4cHLbYkopm/59bL1n90uzqXfDHqqUPmrYlo3zbFF9d2cRxn
kGO93b0VIYcw/Qu6VLKAZ9bIJ4fA3Y+Q+p2j4zOvdX898eVxX4Wpvuv4JyzR7WYtBaH1KSmuYdfR
edwY9Bc4aG4AFGo9bjpMaUNCdhfjamymI15LoPJQHNe9LAxxudwsEcWKlYtanznPe+LoRRilKOzi
x9aZ/6yJWkMhkKtc2mxXAI4pHRPSoqoTm4qTw6EyapEdveqOHMPxIoKYvP+Fbr4LxLGYgmXBvift
sia5lALHRiUUKrvg7otRcfXk6DmDQpKd68HB2bejOmAyqTG6X6VZ3GOGPox385upXpIwBW+w1ex7
KvMa1TUM9Drh1LPTjdjR4OlHHsFErxpAHGAfdrztMVldMg2eAoFgV1pMII65PzxCjnXPf/qYumFF
PXiJIWmnYYDvXWvTLvUiPQNaPFSE2OdvKYKylENLdm7vnmyKjDDGgVzO+os9jiSYBPaDMYpP0wOO
LeK8y6Jpl+7UZsDv3gMtLuUfo5wFEgjSgUWFRLI6/IDONt69OD65/MlWU11iQFgAWbWjkxy38Bho
SP0aBO0FlRRQENbk9RiLRLrBMGWSXIbDtuq8O0WSuicTEgw2GacLatYBVB4a3vgUaBh/FP4wZbkT
hIz7vncrKoPoebKZ33Uc1ohaEebdx07YpaUExT038pC+bP/M0+NPcw/0o6nWZsQwuGrqPrVq+yXB
jswe9dOrIUxG8/N6imKfAUrnixYTQH/GXFZ2Sw2aR/nlMfP2TQMm/DBQQnwucDl9zD17jzHyviGW
75DKGu+qeSHdgmhiXgwpbC612sCQwiSbe+Z6VjHEffFzdnXCL27q5PeX8EnL//peRN3C6B4/BONR
U3xTxgc/K0i2fzCzY/OpKq/R6iBBfrzPIJyRIoMWSJkyKNXq9GCaQV5ylHrwKU/Pgq0g/t6xuewO
KJopybjm8JBg++dMUbKBa6/Zt8WIdQM9K8jvBce7yD5JWJti4NqtnJm/55sY5a/IrVGleKGQ3E58
EvBayp1cIQN8gnEO2PxFNYH96coAIydNEgJk+DWT/QJd/o+/QXGdDVbfSB54HyNjewYr0YIWyrLF
MTXLIPlGJhqg5xhVV0xh0r9Z70USWAVzvcV/9dZpcO1y4tnSbZdhX0GYzvlhOPOJgeJ0dVsO2BH7
/kIwN6pjgAk5nzt2nJ0iuns0NFRlg4om0iePWetNyzwkB9Cq9dgu3XIDc4TJH+A+QofgDrZMPp64
N6OdYTUCYjlyfl5Rhuvz0FkN9QsUNuZ9hhZkGaWyYvWtWZKlewHm2D0U1oHVkRjypvTTdmHwqZ/o
E2EjjZZH+u7QYdAGjLZBwp9fqii5WL/6dEFkuhoC76v5KDj0QHibbBNt7siWgT19DK2jvzjAHZ+I
28U80bvTDqD+6S5MUzj5B3SlKTZw62f7J/VYxphQTLLPUAffPLcHpcKRpwfENO7QxwxpxtoLPGJp
UmeQ7qeKHEWgyHa4CheEx2gALvXQpU0oIWuYsl6AX/6EufARgdEHG7J09Vm5YgO6okE+Gigobn/T
yRjfolbonqfxNjbbMHsonvnp4I2HJk3+EdveUlZgoSdnjSZpQETA8NGhnGFS91bQeltWgl5kG37s
jtdfVG6Ha4NFY4CimLEnaJImjU+JvxkKkxReuvaAR36lEXemfeo2O82lCNkXyBPMieXmb6I5mhb0
XLrjG5WTUuifgfpOEUfRvu8KcXCy7z+4TjcQK5mjliPKvQI5cbsSNsfa4kLoPHZ4Cx5PJYaf+3f+
2wcc+BqRTAn23p21cFpeSq6hdi1/Bka7x8chwHsXCA27LM5P3sWDEtYa8sBz16yak3DPPD6Bz8SU
cT38Lb7S3zOBpxW8kWGn8GEkU9BlEEjP7Cq7decNPJNScuv5zsLXyhA8Ul1XVGe19K5HKYzcSeKA
n4T4xaPu8QN5LBUSrSpGeinUEsBQzUUKgABy7FWOb07a4YIXwKY2WhBBXTLlyB2CZX04/0M+ExDI
oaceXxx3PeTT5TYg9XKWOlxBhCRWN6kwyGhf4qwNwiX2BbJ4Y3v7qLrpyJS1OncAYsUix2NMkYln
5/wc2DEs+gbvz5E1dFIJn8EEzF6Brp3xrve2wb4QZcN4uxkkJtjmBzUhXwc//Y38/k92Fdd/KtZE
ldRr6Ge2r9a85m1svk9C+MDif4+4ty3W5HELXngtkqia8PvIX/xYwK7j3duGlQeGqMFb80e2ACtx
vgHzyqKGkFE8DVZJtx9FsEW+GtVkLub2dLuFekCWCsKvg6EO0nNWOloNhhirdUF0jUmRqz1Iz4PY
Coio2aeGKmuRqE8xaO3mza4nt/9i4WFf6NEarBqD/X128+eRIWf5c0lPuMDgwaZIS/4JOQn3q17q
5yOU7lMAwMo/EHCmy6OZjDGxVp6ROfYSi+rhySpdHVyiYE0npIQVk6SVqaI5yheO1E3fF3uF6thk
Z/BtuIRD8JfASPfib/O6/1rsU6wVTIlSpJn22K4/vIg/VOPEGnRPHwawQ6hlVmyH/pp2ORsIuH81
jthfYgPxlkmFovN0Rh9fjWTPjf9ubaFFO8R2LrwWAOAl7F4lrgRgkPBjdBBCqVeza/sd6J2mTo03
jAsilIGMgxG54J5lfdIiuXWnEh4Xy/oyEG1LbxdFRPWpVMXkg61shn17QXFAylP5jLPh9wws2aMX
8UHu3zDA5ptOzqu2diPZmzULbnElO7g1n1P+MOmn7tGYUjbP4k9996npyY8eRbSClGK6XzA/N/7D
5/NAg0xH3x1y8Tcpv1LTRE3SJlKc8xEb75rT2hyNIL3d94z/6VXKd+01hA/HDv4ocmxCC74PIkCQ
Cnt2mAlxu+VJCYyW9bOk2hk9sTEl4oBFrURHbOB7pYn4CKqZVvgg10IqUCSyvPnU9IbfVVtXIekj
pN0g+RXhz9LzpTGhAqktrwi/WXOt7z41zyH8TtxrU04yavGp4XolifzHbRf3uyQKrluux8y9QiBM
TTTd5J5E4vOnJKT/zEEbYMCrxQg3yrTwVzdD5iiE01F+sXrothEpasb5zGLZgcQb8SwJJHGFf+/J
nnE4YseeDPAmJjuoHlb4T2KXXA1ejrRV63IGxMftAEzcOvifaCqdNznMcDD8ZdzuJFAUYn2Gj92C
9EyKq3cg9mkYP4iUG8n6NeSbMb0BCKaSter6/uHvcO8pUnKLzWwpxLF+CQjzMcLAJ4qx9r+aWZMN
UIOxzEF7/HMTntKuG14DKss9fjSR9odw2G35YPzTy3bhre5kMYxzQQL90l7zfWWkiiLFKV/iCBlf
Wq76Q0cxcvynnuVyt3y9ikJueI6pHPyVcLFQYmG89oZAV8toaXUkMxLENlnikBy604EUFFNSlIP9
9/HeQQCPidN0qc7lecCq9wd7tFuf78qrQToFzU30nuzt4rfpsYbymLdSyma1go/lRNK4Hfyh9Dal
VWRQ5PG2tYBBHSDxZYjwesLZK49bjYD26NXXw/TDi5BIjQdUwmG4bhapQvjMjYgm8Pu/oxiVnV8t
AKfEes56qbbAtdUDjlXQwybYrvf+lhVTNRuQcgzNgtcUSdSej1IcleGMpi+nlS6+xKtmBmiP9j41
1ZKiTUYY4wfQmM9ddw7xoUbOzQa0m4LPDj3NKdtKVO+Hj0qyu410szvgZ5lVofGXk04Ot/tkVgNw
YjnnbNaRLszvrsTPtM7fzs/vMcRSWFMNMiFynwMP+UwZwMa0k3Zgwp7sKtsV8vbOyJyUr6IwiqzM
rlGZhBvFNjZmPA3h4tQCxMoZ7tjgoYHIVrVEiZvQIKjbzgsyyAdVg5IBgruf6uf7vw3U4BHO8v/C
ns8Kpk0EH9O+lckzqTBJQjTd9nGqpEpob4Metj2DlLuK6gf3P4AMvFXTG/fQSdGJdXFR+gqa6Yqu
Lxh5WwxqN4SZcS2L8qQbvkYM2+nRNE8mPCIchW589hCx5IJwX1U8dWYd2C4/JTdMb+IMIm8/rhUx
72Ra607itRziH6/nGa8wN5RGyNBcdeomxqMvjcpuBIvZYe8glkqhMh3tZLR7//QqLhbvkRVvqdDj
oHtcD5kl4Elt4Ar8uWSqFO0k5llCthy5W7CrsF7qMYkGOmjVb3Ko9vdyOP8HUuNhVjFoz2T80DFs
DgsQaG4PqCMZUDqKruKJrGN8zZNTE5K0NRkxB5xu82CxGS2RlznAlsEeE8VToZEW5vMdGuj+VAXz
nV+mwPcLqK/s2HJtB2Zg+wTLJjJ1H1FSkCow+Z0uXjPpxEhLqlyw0GyFoz+o+Gyns8AZgbbqftFH
w2Ur3UMnMK2e/jO+JWPR9ZmNCCG6d2YCz7YTHSrLxvjk1OCV3Dym7N/eoFxSW1CeV3ZjXpEirpM0
Kl+TWx5ldJBlQctHeReDxRG+7V7U5eFlwapaeHKNzzsp6MNyrvS+EVDTVzuiR1zxA1ETrZzbU8Qc
YQjPJ31HldcJ965/CBOQg5IYyDvPnuBfwb+wumxp0wMkOFVBdXm4PUWAlONBKc6UceNs2HrToGMc
S0zVz+7ggjGf2sTSl06izfu7Lblpe7kj0Twi76cEUk7Keechd3VWgXp44xD6qbExzfPP8B47S4d5
8mP6ssr+TEkNqgxz8gDkUp9Trf9hs478I79XMZd0+JBvQuSDF0F2clRdDCE6LjXxVoGrRgRFBnW3
wnK4piLL92C2hze0DX+CHnqOeDwU1J1KEEyw67GGgrGAy+hEpL5oXCyVdiefm8MuPvcy73vWcf16
wV+1W7peT0waa0dftPt0ElcFhn7UyZHxyj5VOwRxTDnnBx2NkvKL/6i3e//DVM8H/k+mdWnuqtbB
rd35lWseupqoPsWzs2qsjWgc/Y/YT2esSXVANA9fhVXeLUeXpSTwGvQczLR6G7nWRkLm9PeSe7du
x9JBpesGkH44lNZFUCGVSXn63745EOmDoulu1msRa9fnQM2RCJq+4kS+4r+NbOCVpPzLoMfb7Ezg
VWH3Bleift1Qx5wXYLVDz+w3xAQ4LgQUT+9jIoWOm/tj6PV1knTU7/hrd8X+zLxNUHokLm+m0NdP
UXw2THTULEF6NOGCYejmPSoPFDNo+9XiTy2U5RM2Zp6GKzS+1PC6AUBHEkOZKA3e0ShNevpB1ou+
QZfM1UU71EU0XvMW5SgGtjNrUwW33flkaRxgSeVz2Fh2Wv2Hl78Tqs4iy75JaJYZfXPH6yy0qMPw
IOTiNSDK+FoONl8ZIp3A9HVGRUzL/6NV5VLzQDgcseN1l4SmfnUrkuvSfZ5SHuPhie+vLy3/ylRC
igZaGBrcvHIDtQdSjENrtI9rWUrkk5axkrqXR4KsuH1f9N2ae/GRo3nx/im8f919W27AYoC/3RqT
AW4s2RMoCJSMgWvqtYVchjyV9skQs/+8l7YVPoijKrm5uqcRYKv/Bi6r7zxCkgDHoUhRK6XL19BI
OX5mpX8CkppZNSES2ozCquI98qwbm/CCDAb9l+FBSIdh2yW92S/APQcQsJ2JKNCxdf/KdbgRp/k0
XwaERmV8V5HvVqLNcStUoB8vfd09OOb/Xlhy5ogoLiW9ivKQvQJ5sXyN4G4iul29/qVHLQVCgNze
S6f4iv3BL3W59rUqk/VFPQdRfy3ZepFOqSeCRkPT88/Job0V0gDuLv8EoHV3s8kKVI8lXar1vGh7
1lX64F8jrn9cCktiayt//SWvQSktR0EEtAziqjzV5+Wi4/tDrAzsXIHzE+Prstcr2EIexa05BXwy
DW0GboTVQg4P5mMjrTY5VOuV87E3BnGyEwhCJLLico86fJTTkbC7YRQ+q5guDovoB3RO7RnvxKwg
u3VRvHQ46JcCHCcMBkpjdhawvj7AFeVslgE2+q0kAxMk3POKWJaS1rWJSS37J6D6+zstHoYekyS+
b2tCTI9G5gTwsHaqL0cFelrpbIND05ZGDvby5/boucDLi9Oodk1AJEhh7R9b1xkJH2FqSPoAjNqm
FIeV5MJW1/rPGy2CQJQKmvkYJYtvv90LAsyrC2X83tM/pCKnq6C4fUiAFHeBpGxOT3ClxrW/2CAx
0gXSvfflTtZuSPD2/V4+P1EHtVSFxM2P4xCwBwhvf502J46lDmYK5udRSP25Je5POO41ZRfwV53H
GvE/RIHh2bhwgl2rf6351CEXZZM7XjJ2S7tvKfwfksGLXFA5M+NhCRzmCv4KjJa8lSDVwIBar7ft
zAUniLUy4soVRc1V2VtWnfL7KDjR6pe4kaPJP7qGo9bNcALoxQrsvQcQH8l+khpFzEKVi1xy4OXd
qh/4+AasI8ANX4I6JufHFL0H/QkP7OEejFX34G9SHP7fRGen3RKjDPP61KdGaE56jFqLYKboRZ0e
EPbvsjhup9/AgE+fgMA0SgXb5UKd40j672dVJjnsPuam8CSMQpNrjYqdsKfVBACxCAR7MF2cqsPm
AFvPAEZ5tM/lTGUc7gAe/iaAxdjNicpp4S+Mow1Ywa0GH15VYAiV6Gsy3dIB1g9FhiXPsHDUpM1s
HSMrYvMF4KgWBYL9SGYddCE8H2PA38cjsALLAAT2oZaCN52utf56gfc9e128LNreh/S/tU7IGtEM
iEE5sLm1af3L3oGJYqBCriM6x/iymg4U03w8s4TQWjh4bdIvTAVqQot5gksUna4goLsdm0pIlU58
M0ye4RiPixzpb72HWxnyY0aqFW6NL8ugNR8c1UHEmuNy9Ii9ORo+Rf9t6a+rxmXtXJ34nI0230sO
WqTeOhBkz8fQVBWx1Q37yotwGnAPtbwx/X2RvMA6cOY2Y9ZAtPzWGTf2okdJcBp56L5wtoMaijO5
/IfWiuA9VcN1nFynpkJPmjMpfaBqIbsyT6x516iPEQGN2PgEJoPcoxbrwPTSfG0g+sRHFFSFm2SK
Qv67bHzV6LIFDKHMPpch16HzMdp5KVRhovziK1Zht671kOn/R2BuUiMmDhZG9HK/IN/c8cUCtCrp
vbEO14Ze4pra4+BFiwB91NXFOpmXUVWx9Vb4G3iCOQvL+zyhkkWDTAK+I5DK0rRO+77ZgqoVFmFE
CjWpexE9voP02S+drycNrlSB67t1eLH6E/SH5AShXCqP52vvL6on62EbMyb4WzZ4n9mGx49H3f8I
4w41dAi51EtqVoelEbaMmkn+IX1R9VHeh4TENj4JPdkpDNYgAN/pSrg5tDwlhJUdLHjmZPbhOeta
H9LN3IAtzsPqQk2p/DMGbqRJQsqUyM0CoUtSu4n6jyAZyNp+gRk2SH/N+6GAb7B+2pNKkFBjNE7v
XiLHS/ARXKdpYC56g0YEsjs01ywauMo0c1iOuq4HYriqOLXb7ajFeSLMFqDfhWr3w2rEaF9+9I5e
MzHKwNKoVHm1ehkTvK1s1I1c0Fr3Qzbj/ckhjrKIiiVMOUurVz/NXw012NyRdlc0UVfEZMDYWyR5
drWr2RHvheaj5SzboCYTEfjaXAsudwZrx864y6TpjBTrfdPgNy47/7wtihC2RKG+mzv34VQD6MBl
QSW+KNzVd/QpIQoNOqmQqQkUY7a2q0dKuhpxk4ShFMVbAEPI94FmaA6T1DhJ/ISAwOaNjoEEfpho
O7H1zndTX+6PNzquimRdWY9Ez1vKF1V/yrrwdmgjsiQc73fwfjZd8R8PlWTOBH9T5+nghsPHierx
gF39cPvDL4/28fvPkr1HaZveLdOzfi4y78xY73Jh3PMlm/NTnst2ZMAM5DOtCDaIAXc5+HS4Mx01
a/RHasa1Rb+Uw6Sdalz/jnK529OdScWgRr3hU1fUBL25nAHe0FGg3HMouq00jwRDt4x08lwG+rnJ
xsFZe+NyxMlhkCHb4CeMUlbP6NJrCAea4mZSMdfayjsWZnhpiGj2NJmXL1KWP4jRvuti3sG7Odjn
s1E6M5+nxslHw1GBo7XgcwdbjWtXAidYZ9bSD8zodiBW5c0vRYzIIo6G1MWSvgcYC9ta6SCYJgjc
leinIKjq9e4zDeCqWriJbIH6CO2JAcUtijaF3HcpBBUcSPn+QekadiCzjNQ9O3rF2Hoc8sBx9whp
aokZCb34Oqcesp8dBhUUIzzv5PSbnanTk0aokEbKM9gr1kInIBZOvqwFb/74mqywlxgITCIt5wrV
104EcqH0sEC7MluZ/IARb4UkM8iKCCGBTJB7erHmdEssmlER3FKk7o7QLnBzzXALTm7/pW7+u0no
WVzbskz9++y8ygWa32comty/DY0vzgPnzpFxIpBuD4N0xGA8PDHqIixVlvIoZrRswuBBfC3D3hoC
uXYvQgIJz3YosFRK8njKDljo1uUxIdeVK0jT9Xc+9VtlGPBa3EFRd4Fw/eceH/Vg36x0iItzl8P6
lRNYoFB78L8eWMLE63NGp+2zMI9laxEcXoMqt3j7RROvOcLG8HSfIBLFOGJsoYx5V9d6sR1bsBTy
QnzZDrQVYfKBSiNvUT4Y/lPZOMbipRDwCLFM1zbLi/N0VF2NtmT2lyqJ+8NRbBPlmrZBAeSH+JtX
EuPXmtNU5rMkiYOkkFFKxLNAL5QnIhkW6VbO5sppGJ0fPWhZkQSiwtHtqiHD2B7dppUN++zpMgwy
I3U6oHs3UCNvZihsVCbyQlVKJUjM5dAyp+8p1otOBowp7zpFitx+lx6eekioFWlERDEXE4l1zmzZ
9D3mrfsT9v98/ewybVzbVofuedLe0hUtR+Cfq6GryEfSW4eidZuUfqdmCaMJt/Jm3arSSwBMNyiZ
CgWklIBg0mfOloc3TcHaiKWyN7zG8IkyGdKvgVDyf3+2HMgpy2BJUfgMB5pF2+2QgvbdrMfw5JfK
KqQhvYgx451J5TKyoITNQlxsxeh6BG9NhpSG784JtqMq3makKhzZM+N0SCfZw7/aVWvztkwrzAu/
OmjE3bB3TALtb72KNmchetmTk/k95zgmI1reoinbYHzAkrqFGOjxr2I6dLHu+doneOzzPr8NtaFG
PDCKH6HzcXxNhxQk7/HBBDtwt5G5BipMbphdYB1ryQwhtU+1mjRH6vlndkfion9QcMbKgT591Ott
/1EG/8wiR/JhMrsqEzQHGnRG8xWOzq0trwmy3u3KZlB6vgi4KevRzeSpvPG89orN90RhM4NEqL2v
RLroKS8F9flliXEWOMAqmuQSc32pQm2sOGsGzz+oahq4PFQ/UQLQkdd/ccVnyEzCR6pDUiB5B/SV
geKZs2ZGWZ5EuCjnf1HZvjhzai7w24onpBDqd9DpZpZKdLZ3aIcWgBeEccgJJtFsH3WmIwwezHB7
um/+xIIBZPHQQpYO+DalOHuPrUBMMBy94EzfpZXsk4GWWNacb02SryZCqL6rbXQ6ar8cYodfebH8
Rn+ggzWkGMPZAwtz5nE4MeoHNulWz9n4c89yPujFCK3T7kYxY05H7kOc7a6Vkek0aY0Dig/iS256
O+XpQbuJOxj4HNxBAadpivnD9aKfshFygLcrwdDvEkvOTRP+ctVFo0wSem+7hi8EsImqwzDMXwyS
HWPMAM9Lru/yBDg43AttNpwRfqGcoc6LtBANjI7sYTQ80RuwUaLj8tKCu/YLRikCEKj0G4PT4XiN
pCSxVUTvRkFizJ9MgfKRZ1YHx0QXMVnU1TgGGxpvCPq0+EDW5HRytrlCGCSAY6tUfKQDy048JRPH
tBm51dc2jzVQ2/xh8DTrRN8GOBRtAEneOzNL6+r04xOInqgMR84MCE9p9fn6TQip7XzpvZSyX/KW
botbrIyFtFB2Ia/DKNBopbrV9r22NFGqeHH6XAT2bxXf4RjDZalsV/lz0c9pH9QB9yU0D6c6l5bp
YZKDp6tfP0dV65uPHhI3B93SfQiTBUTBdgaz5Wcw3tO+Q+PnzfV+rzKvlyq5toUsPxigJXcAAo87
OygD92cqvelX2/dD9EtRLuGBISOySLrYW5xpDekXK53AVwXRYJLVlned58qLwGRx1n3uAHQ9xF7t
PyDcXUivkoe6TZ3zFsCOro+8uqRb5VjUftkBOz0HND821SMNLz6G3DzO9LFVJHllE2zZlsvLRG84
5kFTP0v7CZo3oLYRVw+cq4sC541/2tR25BqZ5/OCKxdPuNK/6wYodg/5eYW5OaA1I+No2rpOqBiy
Jkax+En2t9dxZwLcaVqlaSb9u6zEE+xddHPIg13X3apRhuS6ux/KgSMe874frleVEaA+TO4UP0nR
OuZuomsLkkAl9G/UkmFqbC32HXLL5U5uTaWdqsLuaI+wWSaKOEBNSc5E/RLqLYS+57s7ht0y65Kw
dm+L8dbyl/sHALH91PJQeuv/mkpNjicb1TSCTCCl0JnAiTP6+TwK0MAEJvagZeqfzdBCcQWmTxz6
EEcT9dxR/fC2qJfiTWVyQ32TXyQ07gXGJM71kKMorW+32l9MUAHSkVG4FWud/YO8wy1oQyIT/LJj
utaDBXd6xi7dBVdAzaa5DsWgS5uGMMB3RGBvMei9unrbuwcDsBjdpjniOUy48KofgKDEupxZUGar
Cexd1dnceOk04WCbRwu7WfV+XONd22uIZKPGFLMXtGYpslzLAC2GSKN+/6eeKc7h3t7Rn/nhSgGw
lxaaOSPmpli0uo2UZ/oXok0OyVgpgMvf/P+CTP0LW/4iJ6nrnI/7mB0mpB65vnyw5Sm9TmB1Srmv
OthV5nBH7H6uZHSp08bCzxXx3D8sLSMHwUS/nqGpksRS4TL+rkFSlYKjjYEKgOD9oNo33ogYkwzR
wpZW6IatB3EGeyi7GWSryzd/Xf2Tjg36wRUlNLTzcYnCdWuvwbJifpcCWvYCRQR31heRvag2gl63
5If6FyeHMoTCpTJGA7aQ/PZ0wTasa/VlBYA4cnaf66Jky/QGUgBpb7H91rPZDkfePVW+V3xTDp37
5sV+c5yIvA8JcpoHYrwgZFRkL2wmRt2bu2LzKoMrlH7RYffJP2qj0H3moB8NTLbKBEKbzHfZaihq
qB5jTOY8WHM1saJB+dLRDLw6CwGkhiMujvtDBo9Db6NxtY1PyGkmI4PPpjaaNrrOYKIhVNOofJiz
Pr8wlQMRjwted9J0/iiWQ5EUOGCK8wNffd/mMZvmd+CDiTQr/WG9XMNw3vgPvu0xmZ7lHiDaykRU
uitlSoK4ce+y/GcM5QNgNGXVrlbiejWdQOWRAQ+zdpf3zVJBjaOObXNDqSBlKU/uciRsSC8XRXRI
Rrn2Z00VLC5LnIiVsa3CfjTcx4gcH+/jPBgaf0QVhjtbe47CjWdKLHAFHMfwxYLNdDKIW5qEmSnA
arHaWpYXmOZea+nn3FBUmN2udETson4HYf9A0tqk12LuZ2m3MiAM7cfyLV/BGKggAlwuNqMw2Mfg
TTkrbSMPyVaNTYEoWoMb4ZpDt0XZmcACpFuL6SpYAG3Qnmr2Ux25sPPh7Pv63yMaTj7K7C4wzxR+
TigJW6s0LcI45zpLGUflSJ/Zv7mwJvWkgN9VBqumQ6uIGDqWdvtuFuWxoLojwh14NzhiCyjIld27
SlHU9Ab7PmUfPQqWWo5X+NmSCkxb+7PTYgc3tpyHVOtIAeGFUJ9jgs7KIksy0nEf+gw0QvualGoJ
ZHzck/fj16m98CGw4R6w8k19deaE6x/8jmbldcHYi6CBAhQSKlCabUHd5U9U82nTsNQbShqpSD5R
UeTItIfbM1HZiB1LRGmJCFPBblCNXbPsfiz9h1WUowsD1hVsBkRysCP3jjFCZhuBn0MW0z002k9y
Fl8uMDAV6b+uWeeTBH3dYyGO8SGsezz22YBLNxax40FdOmnPmlv7dK0HyKTnMKpuWvNheWeoSGIU
sAhodqJVotFL+O0cUeoU2sQpnUgLoI8v+0HrE4q25i/JekU/CcRsGjK2smjlX7bPs7w9W5DIVz0Y
gbYdl5cgJ4w6DQ3nt8P2FAqpbgN6KxNbm2NzzCH55HfD6dYJxWow4dIHbJ5h9d35B2Oy4x8f9g/B
E2ibHDhiLVdrcyxtX9ubBQGTGpCiVzeEAVQBPDliE6DQ6mfQMBVYD6QTBDPlwaPY9VcJyl0kgKaE
Gs2ITDLHu52DvQOmkg6EnK3/lfF9ZdbgmqlN8WvuJxw8Gw/Ea+iDVqj3VTGchpQ1cmNFGzbLscjf
iaVGc0KqaOfwB+YLpjB9cKWOpqZDEdSEQyRJIqGikzxqTtCoqWJ94P/u4U58wgug+aGPa97v7XUD
8LG48tb9xbU3r2qupkMDFZt/rw7oQQFm/FvQcZZhkpDWMKDBvnlCMrB+7jvv1+ckiT/cfjA32T/K
VPdQ+uTJGNiwi2mNrvd7X7MvzkvxhjIHhnaQ4lcG+SK0HSXvntJM2+PvzmnAhZJWFc0ZRE24azZI
dQdeu2FkZotwZxZT98t4XpAvvt1blXSF8Ta1O6Pv/jwMd8kjB2EKt0tnuTNT+MJS//RdtGYmjKDK
DbwtTlRyKSXVASGEd4LaYyXbqJON9US8wj9Olpux06en2kf5zphl5l0aewGqEpoWPJc0eDXPMSAh
wy7w6A+4X39phj1oUL8XlnXWe+hLYYRWGkBQH9BYgckxvR7nksfAwtn0HcmlC7IzDVBfJ72QXauG
T9POunDAsAmhmmZz87+GqpNujT8QsfpHd414rZqIaTpubxQxg+m1WHR/PZB661xYsrwJ0ZlpEJ/U
0YirYAzaTk+5QNFCx1FfcLjfyO7KijItW/HCItXx5Whl/kR6LDflh3Kh0GJ7nboNWgQVJGxI6qnd
jqkncF3zJ34M1+6sNZyvs7oWUbtQ2pK4wSAaRiAS+Sx5OzUmvPZBmNgS1F1goI9Zu4T+LIRwZG1+
80YKmi8ha54OKn1QvEoOrJWaDguRyrZZjrEt91D8rnrwyIECZiEV5ll0P3W2reeWlbbJhp+TpzN6
Rg8VKQZihbShm4N1Hsu2H6cWTr37kSf5Sms1axMwGaK4HIidMvFsDNyS3ZrIO6IfG0NBFiUp4y/I
LYz9InhC3ZqmSBn76WpZ6mSbxrvOGHsJRto/LiwioAgGh0e9fSJQQZg/9R9KicLt2PTQWd8RMzfA
qLZonkHVrh8oj9hlNgYHPIUZdwM+5/Q/t1jdTIlUHsKveZtwtKUy6wrag7i02JOMG6ItttETVivs
xL/Ki0Cg4J3VWvrEE9bvUaYpOCH0zCiFHYwHYVr1gu9QGOb7GM1DyjuHahwL096UxIe1sAx65a8O
VKZ0Sf3YeTZQ9cRG22y33mfaavBpRiOBe/kEOpDDbkLQfqKer/vg1DNQ1zDxJtQ1PXope5n4jmAe
WeYyoWYI5Y2uUJ3zTFc8hv+QvgB0YBFSl3iQx+XTFhA5hBmlvUJKi5sd/G4YVrjMXTpzdmmY4e/D
ABRp9G2y2xchH7lKDVthgedz4A02DGqgsJk88L7MByMn+XL7A5853OT2+j5iF6HmeqpYlM+BdXqi
W0pT9fp5XVbKI7aPt+j6UUJ4PFK5vhyADVJTN7taeCT1FKurNNjHdJbcnwnIhF0rNE1Pa1Os6wh/
OcQbIljKaRkGV7+zUPYFS+SAMAmrRraHIipQmFFtDapcizgzR0OIx0qZmg8Na2ysOBJ6an51P/2Z
39qwlyRAm7PZ2Z8IO1aX4pBxQc0GjOuQitoJrqFsnO5pySgcvMlT+cIUDdiUtHYKgw454V5GbWhm
72iML6owZJs/d67nD4/mki02LqxhSKsefOKbNgc9/kq9RXT5qAZCxNw5u2xEqgh4l6IUzTNBS32e
a+8adFwr3XyODLL78XznSTUGmjz4Btz4Rw1jql8tmQiN+A+vIh9bkibcap134+3u9Y38AfA23q2y
RxMqEJuyE6bZsorWqou2nRKP3vV2SA+UM/e3PzWd+0HMFjYDSxovXsRn8VNcXwiBcAMh4CGkTCdM
9b3WjD8oTCGCojvbRHvDCfwc3LWYJ7mbu7audckb4k/iUTzTvpc5jsJkIf30tjNRi2kXkStO577h
O3YB8r9Gpm6i+GzG/wNo3WxNl/on8jbmk7/DKwUKO+JMIs1a55lnBWExH8mSuHUCpZnizrgG99Px
IWmzuAkkN0UWozJWgFGgiUlrJoEf11jDcoyzTVrKEybyMhZpqI0cEc/IE/GGhIDpnK/YUGjjkEui
7xOpLBL/FbQx97Syg/D4ur2VojLuocwnsJmtaowyP+rBkCnhgw0NRGMJEFbcNZwu9x6cLkMqyWLF
nwpOkXDtGOiRVM9Rusw8VSUTz5ZPKZs1MrjIBGNcnnN8ez/4P1A1rwAHIEYFoOCI6aQ8CFkhIF7L
6Ja+bkFTMxLFbqmii3tycBaJKNbFSqB1EdAwGnrxG6C9l4LLVOcpEze2+ldOEU7PcYkcmPaPcw+h
3d3uUKA8n4v4I50JloAPuMij4cw9Kw8YFT5Cd2kMJRNjw5S7fezW+0A1v9RAS/fmxZvVWn8fEakS
IlDAs/xoZUYveqcfm0RB9S7LrPbW58UHQ3go4+nMjcR4esvSk1mf7KQmHUIDjmLWCW6G8SGfqHB1
1qGNl0pbFMuRmuMKlnqmh/b3XG0Z4jM4qP88UzSwvg9hwa4hA4frHuYoz3A/Xex5jvkcj54YRIDr
0eNfjzYDEb2s7e8BbQXt/ccnhZRnEK3jTQOtvToV5iSl/IXHUEnHbA4LKUquDT7V5rheRFOJVfFV
X9E2BdufsfaPFdKtpR8YszkUVDR4oKzAMCrPNEWd+h2Tm01G0A0dhdX114kUM4XfXYHsTwiymkjx
PlvLW5mDE/u5Qd2YsIdp9dIref7j+UNgj8FzHI5XXTl7ttZLUeyGY+OsAXbrUYVq+8yB7Bw3+QUo
Um9+4dTN7pWXyw7tDn4GANyF+vcezxhDTtS0Ri5X6ucrTuwAhXEO66LBnR+TBby26/PaAIk+bu6R
nZ65oRPCySakc/gMIjaZrIBoLUvNkRd4y/CVdjCzk4uHpn2ZrqzS2pj7uIo0J3hLHIhYDBvlf58k
YhrK+gv67z+t+lDE4FuodrA9WCHyFHNna3Al/xXbV79zyV1FeLSJkDtMd9VOEKzJNCiZZ2oY7nnH
QcRkbePx78cj+ctoBb9Or+IoI+m60ST+HMoJ/X5Z/QftkKniaWCj0A/GCA2ZNyQF+dXsaaulK/qa
VDl+xXaXXuSkcxJfId3VhaFHAOXwFwrZFGEJVwBHUaANlCWAHfNweL8t/VLRCtd/GbLc7d3dyPxz
eMnlmBKEi7wuod9w4Bnr/8070urisnD7J6b/ZznX+R/APuEyluWbWnn2eKd9ySwh3+jHYfRLqTDq
UNml0/64PZHq2fkzPPO4wOOmMHjvwrjUMIWEUenpcNdbEFtnYlbdFWlhoGJFEeGgH453fz2LO844
m2MF5qeh7hHj5h55I//LdXKAfsgnbLTdJwSgvRC9ZcseUrxzp6QLG6uyitfW9F+gpLjQyWv8rt4Y
//dKedeBSSEv6HUPgn/Afmf1bp3membuBPZmxRkHBXo2CfeEuaWoO6hsS+8wbYATOVybYwqxGVvu
jjgbbipKrsp4VuRAacEXl7eEPXYF3XQf1V+10GCKpHs9iAMvCk7C6w2I7s94z4BNtyIZvsurV1OU
jCjDrvBgMYY2PERPTYOPflYrD6h/6peNPrZgEtXLiVci3DuvTKDj4VBRVCNLtUJPeJBaKxsRg4lW
mKVQyAswijyRkXQ6CXorpQFO9763lhGn59rVsPrAHAFJOjdvO6XQrMKTM8O00/muA8rhXeJNnGi+
FYjqPXz1GpWYxhYtycr1qppDX6Lt0dpxH1s/MgPJ2Dj/5nciHBxnyV2dOlBaubVmgvBflwTj8Jkg
RKfwBpdMmfc0X0WT/kNBME0AaK/zz8kiFJrzYuCHzcZvghegIQmGWrFVx2lhKUfw9TJnuGSnoCaH
XNgdFQx0knZd4RToWusRzWF5fhkS5iSx1jugqxgXosHoXaSh0U6Rx+DA4YYrplEsPrRxjWHpwpMy
Cx6dq6516HshC8wHh5eXhniaMyDt4CauXXBsEVxyvV4HZ0ZLmDMTdj7mLSG5AACNifqTXZr32gL6
A+acX0+LXsYDFtk5XdAVqvmS2OUhBpWQaq5eYjNOOSoAUYfjLDVhTfnMyZO0l4EPscGq41Ydf80v
PO/VISqNS5fQb8G7KGdFn8iFd6VCQ3yHrl3RkvDJYSdx9oRerlruN1ONzSz8Rs6rGyzssU+WO5uD
gSfCVZpyun7j5lmebCNlqE+qorKCRDlkMm0IvqX22oi8lqek91vTUj74y5tWidGx2pV43pT0So/M
9kcf2E5I+MJ/PGFJ/aVnwfFpY/svQYsx05Q7b84zet/b+Yy1BO3LutXA4S6ibXUmpla/p6I83pyq
HNv8P4FVQtlkXWCtvj8CNS35ZAfLimCdwfx028NGk2UI7qYKw3YlE3FDITC/lIiL+I+JOrlKF72F
hhg6GpkMcaos+XS3Klk6VA+YhgivgS+cgFY5nHdmsBhzWw5RLMDgpa3BceDZbE/lQLmRfi2dXOHM
v/N+CjH88fG/GNuK0KCbAvS4kzspoD/0UkKZuuPd2z342wQcJoMIqUGRvqxNjTzzxs9ZBwqFDdzC
Kpdl5FDk3IZ1OdTgDoFq4Pg2esF+HJJa64gs12SuPUXDnE603mIvoDIGOkZlN49reAVAniJ5falI
UuBWzqNW8Psu4rcLT599K2woawmUn0Rvzvyw7yr7n6DqBhf+vmi2PbXWRrHwG6fpKz1Al7UVUoyl
cytApNPr3cowdPxERq+xzVqRgeUqq04+IlirtKP0Wd1Oi7lLEzoXh1nUK7PAOC3ahS4tmCvH7xnp
Q8Fhf8iJuoNyRETG7/QDSRNTKLS7FRFXxrZ2IeJ5hkfD0nLGp+AwjmcG2GqWJZ4A2hvdH0gfk7VN
o0yWkBRCgraQaB107uQgRBJkHXKJaPKDZZf4hzR5A9pX4qEUXJSvnRJzuqYn3Dyk8IRHnZOi3R+N
/lW9znJ7e8LHv9XMYdCHpPa/yFiV4n5Vjnso/uVBhm9BhP83XYhEExiDLahiWPRC/ROnZeaoCGq7
B37Qj7vcHmJkL8//VvmRj9IdL54FUMjWoWCH1H2GAh4FrjtBblrfJGxgu08YS5UyvwpF5/nU59cU
ADwYdqHSRuV4Z36/yyMRlFxioJw68Q88Eli4NQLV1DtYZ4ZKupYB/p1Sw0+D6p2XTW7tdCqTuMHa
xhoUXct+DeZcNJK4WF957QeJRB+zAL91XgK/SRhot2x1u/7kf0cbPZbX7OjPAOYo7y/bo1IIZ+wZ
gBfWjQ5Xv2Ww6qFN2+GNsAH0EXl7ASzZqsRb78qrojqQZXm9vyRq5H0OmpTHcTUpattNF0v0RyH4
LP5Lx/PFLfLV4Ruj3Ny15U7B3B2giSuSZbgdObyHPeUC/TAGq4gkpAxfjZtata3/rcEXK61youL7
jZOvlu7j7gAlGhiKT/St81woILzuLr2HzukTpJhxwt/uBTNvZQjKjiswkOC/04JZ+Qj+Y8GsbjyV
XyCk8X81ZMP4o2wPs0KWEVYNYz4GqVHSOWuAx5t95WBbuVkmX/pAIXNX236XEy0jV9yke3CYP1ZS
cIJxz9ymiq2xfikXMRmj+EtYZOI2JITQcszOSrPre4qCFQPdwlZ+jrqef50qlMqWR7yE2q7UQe8K
5YLDDZTb9QZzJhXxrJQ7ZJx3HTLwwVMSfcPAcmCQxeZ38R21rpuGNinJfjSL31D3sgRBW19US6KS
Z7pAYjo4NCzNM+2dpP5DZaRracGyUp1rciNc9di2/Nts1F5dZ6kEFBcB2d8+jKSJz0OknY+FTwlu
9pqo5pT9QASY/6wjpNutjqp40r9SwgJGlrqAho9cOrPInxm7C4cawk36uktZCfLMUD+eI87WwqYB
vjmPwlavOPoBGUxZhr85AqknyVa3ORyKGTPI5XPh0ypXYvAnFyoho4nQa8PY8DOM+hvW8cO4bJ5f
mdnAgeqazaYNNjfhJ0kWm0E38UWawZmOCTjrEEmQ0ByXbBsoyxdzUkcdiaa5jRfd2YQ0hgO4fnEz
jTqrBoqhZ/h72RWrYxTtCGYob4d1aV8SMxAvaY5s9kuF+nJ1hUaqMQu4nykPu48NQEMronOfGVDF
Ae5zxzpDnscfp3r1vIqROauAONj5LIlcYZr8MSVrgKBncW73jMYhIX7CqKh4QZSg4FKmfpXJeM7y
EGz6GPgH/UqpOqvHWYr8pNg8351b8KaP+iTEfSAlaiZBgIuZ4ICFLCk1S+aXlNuCAO8yQoeF5Mfm
SRrcBx590NVPy2a09hmh2UsYvXL9CmRgeuMrAFI/RmPuSGIQYSuZsixaDEmJjV4ZyjNzvo8TAQYg
0WdNdtajtLDE4NJ7ZuewBZYhMuO/B1nD9mjpteT/DYOF7pZp32IRzIpFCEOWvtEmp9Qg9ebJ33Tg
VQlbS5FpAUbwxiMuShvLi8KpEJs82d3HwvqLjtaOverb5EquEV0/805xYHfDanSaasCJxhYx0Mqi
7piKSoemco9b6nhbaqEeD/P29z0uKgcmTDzeaailQU/mGRToWkPy48RYgFFhTPzzrQcYLjQsglkx
BhT/AflxTdx8kLmFWSvCBwH7JwFurLNOkJJ1gQ/KMs51XQ6iw9EIBMBq2D2kJRqfmO4XyMjE27bf
99yt/J3OGO8ozwzPhQ4G1NalUD3fBe2cofMKbgNNHEbndmp1Dp3fdvvRvEihbwQrfOI/ELcst29L
PWgPl11ql7IXQ42Ilep97Iya9VyjHi6eh+Q8aYueampwgmiF4UQXplbvwqp3GV1ka2M68ieBfBDY
i6b4ib9Y+SD8exFY7owSS+yFZjZi2UGjnp6+GD9MrXPBFUEVv/V6z7urQM87NlN8bBxcVP0cL/j9
O4OJ1nZ85P8GVuF9QPod0OQifuBGuGWJFX5LA2cxHIxZaiU1YoKFjNejjFgoGZNmZH4dpX91kt+q
QZp/33J6aqEPS06RsJS8d+wrJAyTkpqQzZQbIIj1S4XnG6eS8t7pJKk+3zEZeL4XFzRjhANA0SJP
43nm3KYNo+TzSkVxGq6LoTOwMFTqWEkO+pLIV7aPO/wIHZl301HCrYecTMKNEI5bCrw6T2F8SCdQ
j2Biunpe4xsLpGO1HnTGHbvo2HZPOFLIb0+cPsNlHxR65jnUCXIsT0pQk7CZYUeUAzpaes18KDGv
hHnivF1Konizrls3l+HGXpJN01eTht+VklejGcM3B0MwaRt9ZvTZ6paAZ9agFpLmIjqwJ+pLufw9
kSLfICVMOUJTKQaVdsgig4aAoR7LfRZchl3K+RgFXBShhEUVNtz8BS7nG09VithbTlpuc7O/Hj0N
ODzuENHT7E7jRDCOAVi0BLsPF3cOgk/dw5MGC7DXpIcp1AqgRASuPTk0+JA8n/LnDjmtZzVDnuBS
VpJKSmftT7c/EfNw+0k1mDNLebOTc2k67IcYFIHqHXQBFCWk/0zzJ3fpXknFh7iANxOCT8dbs7FU
ho/sulvy+ThYWhAtS/blN3BBs5AYD3HQLntXdOTHgm9BNMAes2n20k3Shbm98oVcHqLXZjLp0JPH
X7MyPd4fxuJzU+/CWFGYZhdWx2bwMcrbZOpijlH/AIh8dF5TKX5W/zWmdFZjx1F4SZwDoBMVVYR1
nTJpRedE5IfM6zh4Z3sVHZjAogx/mML6TkDtcGQJtBG9CsVu1AWTdsLSaGrYGK8a6e3/27A/kBnB
SLOUEFqZO10rF/WmgCQB3fvubqYYifvkuumsulehDXecjlHC0ViYQDujw0Tkc5orCjG2JS9QoXcd
2Kly2xCPkShVl6CB04o3EgBasr6/TpnWsZkvZBHsyCiOfkli72EMPz8Iz11K0sPSg3bZTHE087ow
SLp8hT8CTli3eln3+j32tsZwvb6oyoEgouCXThkIJGl7jlXdZeKQFsOJMKFF5Izm7xi/SfDgwmOC
wpymtT5VLiwo1UbVzhCCzW/iMdt9N3/fMbJrhH0uJ/ExJUMZcAI5NzZicrKNltwcIrqi+dJMRodd
z0AqCYxHzz63NCrt3KvZeGunLIwHjKoA6S/PgQqdoIM78R6U2zrYF36Y7yIJ5JmxtwPItPODyXUd
V03/VVvMWl8frSaiNuuLAMqZdAudHzg/djoTpzu36Pw4OA26K8pmik+GPn2jTL1bdYCwaXxYXpZz
hJMIv0CLtDe2F0/2FJn8OCTQgOswnXnPstwpO/iRTEW3oLtTTh9ibzeiZA30a0edo+4RgReH7L7/
vGfr7yW/vHEX19yd4464Vp1QKZQRMlj4/P1omL4RkJxZA9fRdpiHSIcmiFNFQaYKZh0BBKvpzREy
ZYdflA1BIVogZ9zoO01cJCuCRdXmbPUJtClYQpmgJakrkBpzqOHYhHwYhK/Wt8Ha2vxBgJDlngzD
Xuhdgp335MES/YDOhYtbSsEXSWUKQMiQCND/g29sDtdUQR5HfmpUhZd8u4RMlEaFQGNtPHrLnWYp
TQDZvvZII8OvznOx0k+7hFgHunoUznrU4WwERU9xMk2LimkS4i1S0GmQGt6dHur35SNwqrlb/uiU
dRtQKjnBwqGEDYZ5RH1yxJJTuXD3pHv+labZUbHa0nR4H8K3KjFd2sOGaZFIdT3D6lj2yyb1X8ME
HRlitZfjRJ1HNT7nw+qZ3gfvErY9sLvR55wHkswpNBhB4lCprTlSLeU6u12eiLP3QKlG6ubXByaJ
+7gi0K3OVkYSWMI+kyrZSSQRTKf3xjBekpjivUc1Rvw7U8Z9bEg37kQvNNoiYsrWJIBR05de18uW
3tO5nYqf0x/VrhRqbmpHBuvsPkzKqylz87gtBosTxhfhvWQg2lCPECROApt8XXwud4XrbG6HAwiM
lLnLAVorg2HBTKnMYAYcs2tEXazteXnTdUw/nIUGxs79ZHqeDcn5Lg672nEsVecZgHRQVjLzMTFJ
YR8GTNxgDjDBbLKZX+NGwSnY39oKDKdNZTzV9bNkWeezKbcJxwm2CmKZLdYudfi5/TtpxSBY+l4B
Hqy3fDTY7BuhlPFTcW4/bvvboUyrkhm6CV4OAiQiFORdJdf0xoXFPnduhrOM0u/OVkiyV0iWdADQ
0wXAD36fNIcY3vB9B3x35oBXgs35OSectDaqaEU71btalp41IQinftXoPYmfffZPkl+FSh7QfB26
CNgyWJfk0xTb0uuWZHNkGpCi1qERm+UzqsNo45HmJ8LZafiiI0UsN20cGHFkBCF5yuubTm4RuOK6
TFHZe9ejgPsGCq7zkcrmC7If5nRlWBQbTqSxoZbULAU23CBH8gGpxP7NI+b6fbdbahA+WlRh6K9O
GYBG+WnXn52g5UAwLCusOEEhPtlQyOwU2RTJMVEpFUznrzZPjatbmCKelPNuIiGu/5MMs7ot6QQU
vL17Q7DCEDSX80BuIMEt+CeUJYJWjq8GfqxLOSG9ZFYwgGm0WBfGTCSrJrLE/daTIR3gnJpF/gMl
qkXsuVlTUjGXHfZ0v2x0SzJosfDFJPAf+b/tGe+NQ6snDz6dPtaDjtdGyx2kjQSw8PzX3Svr/2/r
NXNXFTREoRgcZeWZVAuJkRXUw6HRHHgDcdMR3K5h9HBVXuYJrWob7wd6JbmPqNcZuYY1pa1f0ZVq
dKDmT9kzuY6n0RDydOoqxGFvv8+lZwj3pzm3NRPADFE3HV8nxALzkzxO+/1g1S8gkktbFcPZYcoU
x986HDoL0CHHKcYZDzOilMBh58EUZEUoHX5QgswUGT3Kt73zkMt5pUAZoGLT1Vj+CPZql9trx/oe
+hHnwH4DIu0RzlSga7ByKZaCjPPslXtEOlffSwqfjdRQySwTslEfc402DCKahOVJ2+/SkOfME2Eb
thzJaM0vT1J2n2ATUJqqooyEGPgrpqmwIutVYq2I5PNZRRjBzpGSxQkdrzbWumOl9nw6a6ijcjis
Oxf2GhCruJWvWQ6be0OOpcFBRiW0I2INkeds61zr1NXfEzpYKS7teescypBKYIq7b+aZ9UsYT6St
hHatbpZtgqrJSmP8URxxwALSpSo06LkLvD7tpwIeFAmgeKU0P5QkYW8ssCyrEKQXMIEvkmRl8wfi
Noil1y1dwzcNFYROe5pSTbygTNTx2CWkqhuTEHO+B4FHCOim64TPvYm3MUYT1oTOZdD6SMdZsfPz
fq4MO7IXrdjRoCL+OE5oIHQH/Jif/o3Te3Lx11Bd/JYdC0UsiZx5DgvGE1DNai+7itsjMg2B47eT
VWwN7BnCe7bWq+p7vs7XME7YTq9k7BYOAVgAE4kv7ZCiO2QzdF8PQgda6SHbPFuiLlT2lblZIPQ4
dnM0zKattc2sIWl2OTIsa3bJwGGsz0Mfh16JOi3pvAE1eWYOB4jFyWGWiRF27x/zGSttRToVBvlL
Ql7OeL9U58PYVGVTYKExk2MveqIfkpkqIFB6D3IqXq5jtAptzM+xxB/W/s8fYOX6gCzIOr/HzyPo
kIsLtPg1LbgR/95dQ5wLhMRteqsoWhPQXF8uof+wdaoHLLUeM130/Rq1tnhMJdr25sY73nbXp6Cg
5+no2f5BY0QmjDtyzUXOzkaW9+Vc51zhEmhDPKU902vWoD6NWyGCFC76gm460wZ3p+WG7Fk9IuDt
Bt9W2UDa+DYwOW/Y/JaDU8ScfjS6unawJOft009BbXBZsGB0PA/D9S/+SulmdQOeIg5F6HsHk64I
h7ZIOzBxYPKmHXpsLxgAgp+fCXaTRm09Adeh+ky1cYTSZhr5j6dYwYflfa0XewSj3yb8e9IJkcFF
v8Vp+k+GYBXuJTf7FThlB06Wbh3K7l4NrvfaWC+KwvsY58eG6h9SjyiA5/He5VmPvG9A3qmn/zNq
vmXRacWh8B76QKXYErSAm3EoiRSA2XQhVB2u7y6SoZWGf82QfxmeD0m4tG6ac0diY/Mg1Qf/KrdH
BohBukeRlXf8jne+/g+OWhRGIM8K1fOiWasO6AlYqyuk1s6s/Vn8oofqBlne2z1vhcNyXCsa48Zc
omMURyYLJBlfEcmqmxNYZV9vJexRVQdc7IMDCn3C0vCqKglYPLcbaJwDAIxOnjNegS+lZrgkLaJj
etd+BhZvpkCpJsSi1VX2upjEVb2RIN3l7VqW0ZkaPj5panJqSxxqagXW5JffHrhSNf2zJgNwtCjd
S5RVvj4Z1UfhyBCE7IwcNUDv6gxSD2rgRuJzg5fQ2L27qoHJbSfXa8fIqwLAsvu2cdAkY1gk3tRJ
mbfaTtFdVu2t+edzLiEXH+Gpb0KQXX5gSHUxJ6XxSBB37AN9k9QJldtPJsGMiN+UnkCUNd8GiYTo
9zQBe9T+6//36RVQJRhoThEYlT1z7XbepyAHTTWoA7r+cKbH57/y4sZEvy4w9iF0PaeY54B2gX0i
KadXIpNWRQQdiyP0nHutTFZO8Zp7bO3vNOihS8ZaSq/ux5ZBfTwcXpvLKDbeZQN2WTH39xX6+VKC
If3pSbKrxPm3IesR+u7EVYtEBJTlceaZYJQ7+DhO06SSL6wUzxZdAwyjbz4iAC6EaxJlrqazfOoc
ylV937Kq7giVDx4uraQg0nhydVN8PaMA6ZG6wH6HRD/bruZ5OE8BBCrxRct8lT+g++CBU7dY5FGD
8EXoIImm72KSyWprszxM9d107zkZ73Dy1KrGcs64xlFnxUH6liNVW8EMbEh+AB/CWmSlSkcHqPBU
o/NBrlHCxSYR6pGiK2UE2xtKzqJbZjMaQO72r6hED1QYYTlMYydoi+xwoVqIUMQVKXDuH2yztNGZ
n+5+If5JoZNRVfZ1bbJ8A0tEadpM80TTWhWXyA/O85A/FZWjXPiBalqQup0yZfJNfejrFMqnG36j
mS4Nv48cYz2dmqIcPtHWjLjvYC1N/6VC8GuG5dFfNh5zmIgdWnpSTXVh/XqXTTGYof2R6zYspcjE
BR6j7HKggjFqJtIz4vwQsS0swjb2PvR8CGAZxm8Bgc/tr/97cLDjsazskRceo8eOXae3RQKln5IQ
yEKfatCQS+ca2tmAKfgFCJG8AOsAOroo754qSaN1S/kny6mDjB3KDIbceJVywesHdhHoYp3bFzLo
vDmvJKeCXKG+HzPzvXNKqq9RupH6SZdYGCIa/wYpG54nJAluMMbJRjferKpLZMXlnBjwtVSoA+Qk
bjOePdEnRI70cWBqxtDxhmm9m1YkclI3fb5pa+4vArCfJetGEAShTMHS1S4p0o8eZLc4MLROzDdZ
lHIV4nXHEAvohUjSLcJTBsANyKW3HRTzqTxVSMRubdZVg6bU6I+E/mfAtDnOQiEQIJauOaewsRy8
RpcXcyUAPo3mnnjE+WY0b/8qpzfUeGKHh9fyDa+TrY9bnDWzS8M8aGIy3CrOaxor3X6BPz5y3Hqd
dzX/riPQZXGyhsthsoc6Suru97A2CBzs5ljW2cDA3S0U4X1jrUiDEDxWLkObpy7EyeABBCsf1s9V
A7y8kAaCTwwTlY484pZoqgmeHIkrZZiKhkY/aTM/iizKzGiqEzh9A8yduTDxodsN0EgBC7DwhHwV
j9ZcNlYACeYQCFGo8lYQs7qgHWfpQFIZd6+8HsydZydK2v/okM16/9nvXXHzrVwowKWuUa5tv6iI
PrE+tCH/d/sj0kOOEx5samBYpSGkXJZUNGQRuTaL501xa7isiuy45opfOZgkIXRaULWpfFADwrXO
cuOV3i0SLqFyz31YtkpZNCvSmPvbtlXEQZ43bBWFqPIgmcTN2VOhr+UmwGiSvpvJAgQ3DTz7pSYG
aGMprbQk4pNdgnxay0Zny9aypbGozQwTyt91ski/x0V+uUO3RA/yxUi/DXn2b+ofpR3QLhpHcBJd
CG612KaqUVlr1G4zogsYlK6LgZHS0o4QwFuCueeCEFYFO6n5Ta1jRpPBfIQUT6AhK+5Dm5xKblJ4
OhmcF4Y1ctOmfPMUrZRFNCHw7ZHyiqJCb6Mp36MX/YTSFg4/nFn0ubfvBwtjHzYaak822qXtA+AM
jV1akwL/+TuVBDBrHBzhDpzk2fL97xGyyJx23dqnMeJPCAYAnmMQ2uryDEh8PP0JgYyDzk0IMAmX
yoc2ZRTgjbVTNS9oMk0gnHUkRhuDHPfENW4WETHG3b4rYujyanp1kRYISqDvOj4RsmG4VQr2kd3L
5TbtHCf8hnYNOfWkJ4wjqtzhywADQx5hUO+RU0xqfE2Cvu9ghNs8G8yuwdTgD9cZBVEqa8RkOHRC
EARHxpD5wLayQp00IGGLy2CvKjbUGUnLpgMzSzrVPv4wifTZ3UVBBjjlA5+LSSv+bL0T+qXHBaCj
zt3fimCqZoWn5MeRuVWOu8sAe3BH3i69oOR9p7/jvVZ2eLlbOBp6HL7xa5l1+wMYEajTcYmxgI3V
lPbPkber0TOreDVK20Rxb0Ri/pErTr8tiOlkylHSuqiUh6jr+IEEssHQrMwQSNy9T+rwBqzHtXca
ibXWPXx2IgF92pnfGp7Qz5gy/aZPxnrXdBU+WBqJj5VjNQZJXgJYFqr3YRRhVX6duk265xPoPD/8
CX0DvMrPH1eq1C/Onf5n+udSw3F/eaPq9d20LQWeuSf+qeM5s4hxV6ENDy5Jwnrs/wnNrO8KMTH/
04zdTweudEF/mb59iyHlVbsSFMMfl7mIxYpi7ONFo16fzf+R52ng6rbw31geoKFsC9jegB0Rw/wh
JJV3sbmMlue1DsYEMjN3oJUD8OrgTH9ksDBlr59IbI2fjMPA/1SRoOTH2q2HC6VdYH8Ataa6pAQE
kq0QikqjsPkucq888bfgkaAxJWnJ2LyaEzx/CkBsxFE6Sp8V2+CdEICR+7mFJ2KhndtVFqZO+2NW
cdiHUyo13KRYjlsJvNB+z6TrIHsmwl68zRWBdBIJavRTIm4P2xcwk7HTVhZ5i7F7z+C4nJe5cBo3
mAwMw11BliZ5cOkPD/Q7LUUg+2Fac1kCZK4gA38YX+9JLhfjsUXr8GiarnxfIAbNaEmRQOL+tnrH
9QSHU4oEn6YpVOvUPu/nkC0sppC+IImvVv7H6IuzIrlVI7GDsRyVbFoO0ASAfxXmA+URwq0sbGvs
ZSArMiL9ITuhDLPoDCfKQfkNTzOyv256mPRU5yKh5lxI68k0HZko13QoOsJw6azam+6bl7oZrOmO
8ZXr07S7mfaryJcK0GJiN2aG2MbKRkIvzcbx8txDk2HfdWZnrd3vyK4BAjtWn2wkyvbtRFJTWL03
9RaMP2ZMc4jG4IXsXGMdoXkdYAVxOXHTR+Uxj0ygacGBfMsISR3Npu8NkcvIajuwSeEgrv8xLvU6
5wh4eYFaEyYqWdPvpTCop/7Rl+1jLBpwfK+OhftXmYdHav+UZTuAkCpYZZCB4JHFTg1Zl/UxIRhd
P4PRhb116zsDwqGMweJRCPFSXYbMGJoFw2t9UqyJhEefQmDUKpT2qGkGS7mgTj9yceB0fZCLdcw5
R4xN6itg4vQwztJq9tTyHHW3SO8WMjDa8lQr6aoex6XVFvTJfdH8mdZA9nRDR2byRPRzEr9449XN
9BpKdovk1/yl5YbwkB/yXZX0QO2Z1JD7DwNdMfXXyi+2xgC0W+4ODqSCd0eM2OY5vvg7H6f5dDbv
kk0sT0c6jejTVdJErFnN/0lIP85Ez1ln8Bi5QF4A3WfiY5ZGojyZNrDMYuTA6w3mbmT2yPgYSbD9
NOsgDbUwvOtdU0ArqiDaOU3BjRQLc79oJ9N3SZ0Tk2tLAl24RmvbwJecXn9KuR0fIETQAIV9yfvB
ppJwrMVHi2HGuJ/AHlsujLlNDdkvUl1WZ1enZOGHrNV8RiPnwUruRWSPgKLmgWDdIH+RP1euoDtp
Ix/tebMsn6LDJGXKDMb2ldsUGwETQ4oNGIYVIvqncrlNh/MV5jj/OH+fVvmO8H1kQ3BBRrYCZxAa
sDT1eiuSv3anpa5fASzzcu+K45a5S8zBFUHtKJk6Duvz/QelFC0ipMCrjXrL/xqB2B8jEo3vEduF
zSr1xqaW++69HZ9Sjjq6dX6DgVIOkpMcbkjjWCPZolDH7YY8Xx3TAoeLBZNW0WRqg7A8S3F4USFJ
N/4Yycp27D508JK7VW+eY/6P+nxCyt3olVPBQIcop6rA0Um0X07tD9rVR7RB1MzzvxSDyi3gIiub
gqIRAhqo7MRZT9QdatnsmaAWyyaBr2pXsj69Pg1KG66n6KvgG6kk/TE1udJsaSChBrU6ySkNibHI
j8t7JIeAyDJv6r7586xBZ47ZjrL/4YnYCmFp4NIgdpVjU8ZSiRCAMZe9fIPJgA6MCIj9gsKySM/h
gtNDekHcKhXpU/sliu+eqylH+9CM/cga/wFbCPW2pbr9mK/EaiUDNAD1MOfgnKrU2Yy+++UeNL8s
Sjr/oRt/DhSYB/3YoimPG1wpsBpwbK/cv9IlUvvGKo3qG8a3m4y+9t0/pXGgycbQZHQNjntDcBzj
7THS2KMW6wjhS/1KiDKlf6ZAay/w5bQljBtnwuG6bOhOw+GlH4gZpzgRX2/4K1rW2C58yKs1Av02
6Bt8lQ5iumIsl/4S1xI21VB3BhPqyvhuuFRP+rYxT6Wd3wPhtofta4wvK3I775349mUiz7Crms+Y
6InaHtuuyfBnR6SqHa/JycXTEJnV92w7cq9yZUpY6KWSgzxg2oUjcirzQ1FGC9EbjkX5nng6g4jN
nJcXBA8lagCqnNVcVVF+kkqHUxeWi2nKo5fWPPx+85vbwsJoyV9L0fHF2jGFUh/3kj/a34EleXaN
sQoMkxN0odUd1r1aZOd6R5kvMRDki50fA2oVPypSS7cfBZrEGxqp1IM2YVGHl/0haeLG1vl4hSs2
I0pwUlB2og6UuDUXAkohUKmdbb0IChEsvH63qFs59TrpcBt2RtOwKbX87MwIgFVqZIzPUalRlxMB
43oFl/MJ1801Hccb2eJxL2O+0MHmoJKJ3kLfgs45Pfql9BvjA94GqDzczzi5r8wA38D3wm4F9T7Z
825K6/Z/QTLLRYIQItRDB2dgL1Vl+qEDIhzuDCEGr7vPKCqHGj3g9h62gdF5vz1cMYwAzteNVO59
iQfAZM7yWDejd0+i4SU/v6gmLJ5SefiJO4k8850G5miH7x8rr1/zklLPOWBHiQdi7yjTLraVthal
avvjG/uHJ6ddVIVnt+11JdWgNOjhXr1dBMVV/nRRptYe6BHrJIpdoUbyAa/FMBUJUh1ieYn2AdWz
yFUahsczwlMiglxyuVmbMTEpY2HSEBd9/NDixtMqtxL3yh9WtN515xolutI4YTUho8kgrCLNNWi+
CKwf23BKsTsIURjkLf9aTFSKH0E0nTQA+xyh5CqH4egjBMI5i3IX7o0k0Wlk/xTkGxaqDnRx3/AD
IT7P3jwKeOXdrZwV9yN5Q5+t5gpcLK7va5uprDkIzl37Okcl1SfSJT/V4cYkklQRkIzmlbYiqN7A
InIX8hCwulN6qiwVCwiDDubQvRNfZzbTHDFkJV3R6u/4oM0l7z6i6TfX38iNmeqAkL43pvdPkMiI
x+zfEVeWPoUJoGXr/LxWpy5S+n+FcCT3+cMb7IzXHNOOoePdC7QKGq8jpHXlB7LhQOjWSK1QrnCe
i/Qt8W+7IilUJ8nU8MiGT2kNt8W7SaS9+T7UAMMRTKpXtN+xN4HQgztk75XVQfNV52C9X6nPpVcq
IXaEfaH/JdqYymtK8xmy0YJzA9H2YRhZzHEMaS5hhqkyBrhmK/H1VfHKTOSRgmHNsHSpKMpsYhq+
Ni80/6Be4OtVC+174GOR8fJqAstRyBrQbLU6d57E5Je5sbySQ/7UfknKEBYQ/8P8e1YN8NPP6v43
v1kO6PiKfGKU3EuGkSxCICmN1hfeoP8c4A4TchUHYmnd6uJKxtWa/4zrSwUIMC17Nu3TiW5d+Ez9
WTXThmMIBaZ+ev9kNI2wgER6jwEGT6CSJ9zLrHrlrRzr1UHDaudzU+YV5ckjdNsHH/4f5uGfdNSP
1bonl6qFu1+ozg76sa3ks5UzQo7QU3z2awBEjP/E8j1Gd2Ltl3OUBjirH/tktA03z6CzuYo2OnhX
8rFlFBKfQHGVhPNsEa2ccsmdDFjEnodsTvHYetXUwIEXA69owAnbbsvBJRPX/T510RkQcy1YGJuR
CetgqCLM/j9WGJyobEmGc4gBjMPc/7hWxQpOOXHsGiH4zizJ157yFQzIGz6sEuAVTPQdo51r/4Yn
sH1rzDpuVRlZLQWngSHq2BJinT2dUVgaE1czo1h0m/gmA0io+ldm/zN1fkJkTWuLG9I8iS/qHqb4
661CIslv7Ut7aImAymlxjQIVglVMTMTFCWF0gNMv3WjCzItzIiyNDtCo/q4XD2UZdoL8UcmaMrx1
FILNuycFl/Ht74K0Hy/CG2r6ZXpl/109hfRBF1tChRXAN+reFyZTUt5zATb0r12xTNOK3pbk6v2t
giehSvtMqGshlSS/M99fAvfqbsjAMm2NtJeZH4ic9xTdWcH0gQBktDkyhR6yP07WWyxz9MK9lzpR
oVC6h4YPyw5qOo0vwhA9Au4kmFDP8zMGfUCDpgi6Y2pgj2fuIxvyNkbzvrIIhiD7gyN5sadc0vuJ
BV2wN0AKqT0URLVNW1fexdVHidQpe2AWnYTyjrCtyz81AGib8l0y0f/7cSgWlhmxzydDqBT5+Lc6
QKWJPfB5Y9f5I92jdFMqpBfH0JAs80q/nyCJ4YtsS5Urb+HfG83yyjAlP+didDxTJoYAHMGeCdtW
PtLFFV9mdwoKUt1U6S2gayISPHQhMPcxx/M0dez6L/YJ5psHW8G5TSGaqV2gWWofZetCZxVa/aNw
5aJEr0ciGgZqDFSeSV5OIRLaCO/PsXIw8FPRToumcD5EtajwTbF/NNdjRpRSVYvcxhbkCehrkwUB
sMZ4zUZ/b51ANcmEA5fyLrwdmfH2Gg93aGb/i5n1Y9qDbwr1usja0JQEa9GZ4yWTsYWRTe217K5q
+e1i2Le0tf3xisscDan2A3GaevNd2dctsGwPDbLgVp/FxzhhBHWj8TRHJQtYxnGaI7FI+AyG2rj0
iAHlFTYElnaBBPkVFCMoKVoWf0t/AXMNzkVWllnQ7Pf4L72TMU57CbRVzYglHj5QakYC3TMO36lR
8XjNQ4VgwoZMYsmUGFb685pHHjC8iQaa5ogwWXDfwbRmY1iorDOeQg6ZeSSmaaJjrcyRZCfSLxY6
1DGFjbT9uGwIJAj17/g+ubsac4+U+KREfNAEl99qnbRfnjhLonFjNXfqpjuNqfs59NYGDqPCRmH5
GXeSw6i9uJZoZqiGvMn1Ryi8ucA/ave5MyjqyjTc7qlFO/az4m6sz/gaZuhJilHZFmzqPVgHliBS
kunz2Q8kQzY9PFjMlSlCfMecJlVB7SkAz1ohd+MlPlw2cwBYRcXCOvXhw1gARYs4CxPNsoWAUUQk
5hDrOAEyMbMhAbYPL/bmDcb4nbM5qpsFe+NWPaFZU+R01nQpU48nCdJo8u5wJs8RwCzYc0rhx7pC
uUIWIJlThewUwhBUWVFe5jbJhFTr2e2MY0OwS72/A9bUR7fFbfOFRY4pExko+gECmBU//jt+Q3ec
eMxa9BGmuq1sjm2Le+/ivOQcIylP1x3+MdntEWk7edYwGSipx7fiGX59WBRx+p/D9jKdHISwyukH
KG2Fxaaj+vlgIgmFLVgYf5KuOU9NMMs5n/pj0zx0/Ax/xGex2kNhRe/8Gxezrm90aTM+/y25mxLJ
e2BkUuvw9Tfp1MvHsr66PZ1YX8KxWWDlj5MDc9n7rCKVWS7sPNSLAEnDKyI2ZyudVDWMAD+6bZ/R
9BCpJ4OeYVMEMGvvw4WbQPibwZvW+tDlawQiCQPf8UQYNFG8NaxbGTI4N8b3vSBN58GEmr4Xw2nP
QlwFbE8SrgZBmTsf8tyUnAqpJxSj9YeUz+QBzkeqxKIs4b/GQx4G4nzoJpUcKnsqdNkMUITJthG4
CTw6jC4GJDDZTy2+m9nS0JR2ceyYomRqO6/eH3AdI5T5Tz40lrHc4wSWyG6z8F1qkKSQU9P2jGqx
gXqbnr1vUxxCzIEsfLq7+BJSiwn2rmQgUkRjKNSM9hhVzFWnZqv4JcUu9fTjWH3eEfEJGzTw7h6v
lQAqUjnUjcPfJM0UaL1GwnO84aTLg4bg7Rvrdbn40gbHeFSK15kydejhb+Ds3zy16+00BHqzcFwL
ojsDrd7dSNHpYDUj41DkpDt27mHRBlGmoVoadZajQM+fWQUDHJXS6BT24k2HgACf68fm7pj1YwNg
qqQ7KtofIGCxYzrwouiRkvrYQXHzmuL4E7VP5Yer7ow6YLwdwvIrn1qj3b8HW8eT1fh4SrhGRPeG
yMOAIlBrjHaBzhRc4/45HJnlFoA+X5p7/nrlleOAMsfLW57jNCRXGW9SE3HznODJ6l8MSXDwoiQi
inqleGU1WpFKgrC55F4PUOrKDNN12BbD0pYes3fOeAI+hAOB+xdKcvzfiu/BqBdgqQ8xiBvOTFHd
gijsmdP+Lp9Hf/c4a7cO61IVVvtjQ2puSb3b6WHQTkKMa/rquogv482DGEYiK/aACiCFrgZEUfiP
8gs6Wmz2DFFIf0X/ykFECTORzxbtBtncriEY8KRLS9+XRplrZnd2toh4SoHTUqAW6/nFmHmsXSYM
8hfIefOzZst6lIMs3ZDUeiMq8vn5BWQtG3v+celNRbShDlswg7x2k7lGaLSKsJWiOidDO2Et6bzy
i33rkRj+e3Gt5eJXVVwdp6Wh52a7mASuJVzmLpk1vrjN0rJFqTtjZ19OnbazbCfaUlw70hhw4Dw1
oBfTwY2Dq6iS+gFcct3MtSTj1wSCrZ9M9y2s+1oX7hgPWSDC2PWftITa1wY8rdHzwf2UU7wvlO/t
JrMljFx/IRLoECc/SJSAIBHrxA8T7RFHXK4PN1LxGnbfHq3RZbtg3xcod9sZZLK1U3fcmPQqSwFC
pI62RrKh+5j539NWdu/5mMJCpZyN5DXhw1EoLgzhS6vDa02NmyAJRqyiiV4Y7Ya2oGks+yfxt935
nr6pD+5gIOXES8iT33BSA+JCTgczQYhUyImPZjFG6g1/EHBVvRfp+5oQEzibi1rs5c25E1BNUvIJ
yX/V7ZNvsit3wQmzcPyznLBXBPYW0TEJ/C5FIiAwSr4zZZbXE3hDfXwGUgxWuoyYnnCCByOtH+Cj
ZK+PjdAGgBAaG0m1+QYXK94S7A+xv/9t+tDpRW0QICJooqp3KTZIuO6XFdW8UscyCtyiwh+TUpxr
ipoGGoicQIsbBnSh9/wSQsBT7u2Yy8GXvXtQzic6QoHDkXy0OqBHvKCSKrCLv181jjzE525PGowJ
Z55MO+YMZ7tex9VRXGQ23XXEGUW2pKhCb6XYSw5f3JutJgzCC04kQp7mdwGOQA5eDi6fBCF+N1d8
GkJJzgjy65E+U4HUzhuW1RTxEH2m9Y2s++SHK7YwYYly4swL6BTmoC4n0JMT8f/a9m5SryqP1RQ3
ygMxuR4HBP/t+lK8/gO1Xn3dllkDD4TydrmX0y/dLflpm/Q0fHlVYBv+1VSytNDg1kKGjK4pS4DA
qUbTQqKmuZROlpI6DzJ4nfR4P8lI/3kB3Rm0QCUkelEiuFu+foggQJvjhBaodmzLzOF3piM4K08l
HmvoZF0O5ZpxRdeFoNB7ZV/KDbZXw7VX7m1kUR1uaVK3b/iiiWrFVVYIZsKg5N2ImZDjJ55MPwab
EdFYuKf4xh4VndkkHZDWutX/Omw1Ce9GR/qG7LRHMQe3QiBPpX21IOtvSf+PFUua1qM8Y8gveUYj
Qq5lawEKG8Qoea57UmTkj/ufhT3EO6MN2g3rd8ud4pY/YodoCQciBgZWWFS9Xut0/MBVfxBSFtZK
BBhxjEUNGrejqGYFenjhKAcsmV8McMA43Qi1SokEpB6d9SiyM21Yp027eiA4wQNclL2+cUguz+Xl
4mPevRfQgOG+/9lwxhm6erH1AKCJtidgO3Pl7RzexaoDvfDunAEWsXbZUMBzRjSGsMBfEDWvaKW4
x+fFECoyTVm/9dCKN8GWW/2GjrYzF24XNZyxfthl8Q7ac+j+/t25KbA/8Dkohf7zL89X5eXJquJx
hqCTyP2UCeiWfIJdspS/BGjFUI+eWfG+AiElyvGu57ogHnQ/6OMjopmTPytqhZyMicxZrIw4GOgX
1tchQtOnYc6cLe78auDJshdG6LnD/OmR7hBD7upBOjCqZMkkpgoBOMBVqW6emzYovRaHpWRUAewQ
by6V3z0KCdVDPGaZvf3OqsmzWV/cLh4AfXxIC7Psx3+oQ58s1pmL0lIFgf2KWhvDI/NPEf/U9ogl
56XVDsK5S+oHOuS5HK3gT30ri2FsBnyHKMseqHC/mHnBcS/fVDCejb8M9lB5WoM4/uEyBITthC7G
5sq5DkCyIsRJpKAOplt2O3jdBjrYY3iYMgwfszBs+MB0/IA42mUPShdIPYMKOVhTjnXgEERuzyuj
moNi2b5ZINNUwZhhbpkKQa9wVQQLn9W89b8aUz0Sa36e8q1DL/QZDrAonK3fU6+gglmwq8Y75Lor
XBrtmEmW8x40DyhTkwM5k/2MRxJs4XxEfMSaZOX3Oi2d/wIKwDAQ/l6RnRjmUNu2xSsBVYwZVGxi
iOw3PjRS4KBpsV66uSmiFwJ6dOIBinn//x7QQ/WYlznbp0CIZfF7ctvkK+djYucNsC/PVjH6oqYj
XRwGnlrHlnQ49C1kMmtDuY/bowyJfGZCPkKdLWCBHvKemoZA85w2FsEQgBDtbOeFXactdznFdJJJ
krs39+e69OaONojGqvnqQnIBWbCi+pmdT2Bui8D3FGK9sqcFSAyQxyusbJbTYUTILKVnOwVmMnQG
ImvreaH2r9Z4um1km5nAum18c1GB80XU0g8/d3zknWEtlZsFJsUdZXkWTAxs9TxTyT/o4otrQDYb
9Shqq0TJJHWAxtnzpMICW0bIyJ9KoagodB9rsMyW7aAkvQ43xpYEO3vQP/DI7xeZdqdtyn+oOLh+
h3wFOAz29S0I4VXcwbqXiL0QpJnSjqZsfePFgfa/KNSkPEINH1YQrH0IaJoe9QUWcWahRkQRe9mO
h1N3qBuAM80gr2LSK/C/6w7Lw2ZfOSrjDaiw1UuN2OUOTeWBhHXOuETzN2blMRArjAuIwSa8oPXj
u2cDZkWf+FH2NUphCn40embZ2XSg/HBMqKA6anmo5Q22eLDI75UihI0I3i640OAtZ6EJofo/iUsN
63KrcyDJN/t0DujmJjQ5IyEvUvrfNvzxIujLbpcWHLGgISK94Pna7matcevNxHqWGpDjiZFe43gi
7de8WNz4ZrzUQEhN+zBbxFglX+DSvc5TbZkzPBgohjmdyGVsOZpiTgr6gRsqBYvIhLTM9j1JeObP
s5N9MVnV4Jy0i40GOw7RWlnvNTL4zRqNg27rkMJt5tP5FXoutiZTNfWnpMweLjOg+14nWKpnUhuI
YBg+mvdNoMW2keuDQ7tMKOfOvhq0utxLOyJfKAvHv6VPevxZ1zc2wZ9KJifg0D+XFxRNcHIfuRoT
0pCUytha2wu9xqtTU8wHoLUx1/IXP37SKd472d16Acx0mc4BFGyB1ep/4EIEmz7ibhgKHqgNV+Iz
SPQ4WSZJLGSn/wvXdf/fy7KK12LLWV6if5ny5Y8QUGgtHJlPHCCrCsTOvsn+kNiF8547h9H0t0ha
6MPHJb+A2fpQzSx2fGd4q5atPEo/gaGF6F+nHQAB38CS886Aq1HaPE2mRY7sSQhbrtqMtBEY3Wec
gawzrW9yA/Cw8Oypw/EED5ZEfNtrh++WJjXMslgnB1x8/IxB6AP8KGhe7T5w0jM2cfZwhpndHm3p
4nbWnM9scxMh+qc7+cbFnbzwqREXvq8Kir5n8olDDzYel/qsCbuUevHmj5qyAaRtw2KAJ4o1iavj
3ckUfcGRFyipsNL3M6mEqM/u2YPow0NJkGQPBZGP9G4SkQ4BeMZnVRZfNLoxeewBB4skMy1SUw5i
pm4Ki2kRgEgAJk3rI8hzvnobglIcNsVaoXohvimhsGHiRqKNA/SxYc7kKa8yNJpd7y5PdpwyVZ8E
x0itkg2JjGQidg0z+8TGHL2M1c+rzFaxxPYGXv2U5xgOczj1lZFX9QTwiXiv8v6/Q8ifN7R5Vn71
L9H5ANn4MNlcgek1QNtS5bHL9ZZSBBZPXkl7x2p6mTFCsPeJ89bzl5EKOSN/yhxhYjjjFvIwKY35
4Ln61I+cfMZpve7DLY1vhLAPFVweHvKxxrSyV+iLD3EM10afSgaOyU8JAwopq7q5IbFmXTCAUiFQ
/AZz6tIP5Zpz3h27V9/Ac9O2d59MGSYz3Fd5C8OlFsGcoT9Kme5nXH+Ip/QddM5kQtWtD64BjBRZ
UYusOUu+35gdt57D9BPkhZ08n1wadGutuEg9igDjQzIZsF/b91/8+vKaAf9Gbtohv/GA+RztoiOI
wegL48TOhZ4OMkqU4uZ8dUVuCoRPUx36F6mFUbQWiz/LbNzSBtJS/M+S6LqWce5bleVJuC1oczQ4
pKPJ/BSTJpdW1NsaBGIWhFB9sEhcKgTcbeild7ftvPC5GeGH8LW881mt/UjREKB6EGFlh7HFOs/f
lQJxNa6QXybNBpYiPiYKhDDOHPnZq4GisaaGIwli5NdPiUBRimFvG/y5BcZ2761CI4XqyQ/WPGMa
hgFATq7TvW6G9ZVKjajce6GMQDjJTQyA+iydEJaU8gW/SaNqsZ667rkwK2ZT9MDytRN8gtgBc0eg
rITKp7GHJSqOsStofG51ZWBtKeGUy69alPBOdtVx1NDvbH6X4wCksmamJBAbzIpRKJxs15sOZ/hj
9d2opZEwmRsWosDYXQji9nL8S9/RCsn9LnRQ869X25M6QYhUWCl5PXK7RKjobwRLJIIWelKqbr87
ajzuJocbal8iKb6aZDL2UQZrlLFuwBb/qMmmHmD9KTu+uWCwXKauXVUKqKjINKEvVL8ZpvjegJrh
pgj9zGz55mB01YQ0E/Xo2VD3XMzAGghOQNdK/K1QKmya0l+zSVUq0lvGebE0Ebx+ocxQ/+6uyzxG
OHnDB+nzUK61QAgE/vga4DLqN4vQLt1zkxG/9AcM0j/P/9Eg7aRs1T7yUNN81CV1fHNT1e9AekEB
v1IAdhb5DuZ1+2NbfDChg+4q4SKMQT/irA2RIeYe7nAzzT0xi9zBe87r1+/ayR0cHTY3k5UOD7/5
vok2so8XIDlJkuU4tIB+zNFgRD3yr7z7SdTEaPStsEpd2mR0cc+ZL7nA7CgTyte59wOqtF/G/ARp
Hj7vV0kfF0y7OSxR0hzYVhUb6IVZrVU2WrAvYld/0JQVvztX9OaQvAraD7rKohNxDbPROHHXerI7
xiuzpO54QDKaoor+sG1srRehMMDhdMqPowk8NGiHJI3mxzxxnhYuGB02OdUccY1L2npzm0WtqSPL
k3/ZjBJph8USgkH989yVrUWl33Wb3panURdvKUVU+gRno1XSVSoehTh69Zgao0dBoMTI96xwP39R
+WeYaGRoi8HD2lFoUG/juMV91kpJf3KDEhUe1aWCOQt4w5xK8TvO7PARo10encoFYeHf0FXHly8H
Dpzbq+f18gNsdUbbM2bv+BlNjYZu7B7cPKhfoPeWRlxW+E3JWW4gqstQw/VsIPNx4nL0AWxUGkIE
JAsJvc/U+pYf7kE/I3hKBbGgh7SNvJqd3wCmvwlJcG56MKY7fF9cu/q5hxfAqi+Cv84/PJfoq/bI
x/ECctKxUxPvh7KUA0VcqCji1bwIQTODudDZxg5/AwsaeSpeD8MWOwtRNqKzmHnxuTtzlxUMkN9Z
l2gR8XpH/7/PT5FOFSSTtD192TtY7Q67GN7pe5SkMM2urm1uJZ3Zbj7quv59N28LDtsxqroCAx0b
5PF7DF6P+y5hRdvL8oWWs+HkD6D7khaWfsqZ3RJL3OwA3B7tXP2Ur+f1r7wLjCcWVx0nlUg101Hk
3UJyrFNiBKvN2VA0vYwn7U9/SPBMAF0wiLeF/OtZ2qy/78eHy1rLar4GsSAPGGH6Ox70UXnTwGXn
/DWmql7ym5WbhgBIOYiiF0yRZzUgbr0baL8eyHBSwg3roiFDeS8nmOCMuQThDJ4PAAsxLsf/1pAm
v/go9p+V5P+2ZPu07njA41fh+tONHRON15bNHZ6HWu3wMnLb17414SisdI62vH97pXfwS/e99dYg
7iJEDH2zuLZjW105/QuxaFX5Z0JLVanTpAyXFybvPSt353gz8WwIr8AABAy3VCmX44ZDShnXiBZs
5YGsaq4xuDMamGwQQxhMMCw+ScWBZeEtr3/QvCf83p9PGURb3vDxI9GY8hi+EtjaYV5OeTlxGNej
w2L6NB2fuz/KN5KX+KlzxNalXfGAgrLjPXEjD2e8a1Fw8AVKE8EVEDl9rycRR8uOdCMbn4gFLGpL
u9hDBmlCLoiYWUplxiu/k5fSblYUYvXhkQwKc7ulI1Y17zZNx+acbGUcdQU6+G51tJVhU29wXOAH
sXcXTzBSs4XU8DsI+p9nrP5BaallMoVZa3cjV6sDoCqt2h0EbQClq9uLq3M/zTdwlszxmi8YhHQ9
0waeeAReRp9+3+8NYvFKLrhKMzmY1fzUcNBTflefRGUs354+fuQf0tx1hIjze7v+mo54ueEcpcIs
oNusxpHA+zYuexfHJOZLr13ApGx/+A/u00rmPb97GbiOl33iYF+YT1EAZTLe74ZhG8o+OakZYAWP
yR38lw1s6gIQ4hRh/R3AtONKeY9eFAD7RXvrJH3WJu3rPPnNQ+VBuDEop1XH2Nm5QnHZAIQAvFLB
O1o7yF0iSrLdbgPgi1kSF9ArDYm7onlbwL0HKrK4F3AEQK/z9dM/OJNkXTaz2msn71+zTyuGU05d
GV2JxxzCk3xU5BNo/OmU+6lldfgpjNw5MSuNXF45A4AzM1ZX0FvFfq7IwlNNI+3Arej1UOxc+PEB
0ApGvN0qoKcF2RePO4CnW2BLJNb0fTuXvdX9++I9SUVISFm1ktymyqiX4DwMyv4k+u8p0PehWi8y
zddQ7jYpp5s1vt+gecaGy0doR+p8gohlydynlpPrCGx9I+t5xXe9ks54xpQ64uUGWer76D6+9ZFE
mA+4kvUEnfmbdRvjyAeeANZlwv2obif5JaAOFC9FB+hXdLEBgwSN5ppqOOHIAp+lOKiUGmFtCSNX
ntneNVUfB11Ia5xWgdBCuPK7ds5PUv10VegvqRkvWJMQnYr2RPiw9DRS4R4hjQhtKjI6PCzNIKcG
i45rMTl5mqASgBInpWVonIXJcnCz+tfu2X/zk6WIwnwiBx0U7tit6Whl9DuKk74soS9L68jgZOa9
F2XkXAKPBKfCB8Jb6i+V86kNeMMAJs3ivfoYbIZPPuctEAwjjJ1bgfPB6R2hb3YMeaNoyocBU3nJ
LrMc0Au4yMeXOoDUtpB2AZ7XW9y7mVeul6QztMsdQNrqd+meBrW5DJP+OfOYbnjwm3ZejrAjSzJy
7xL6UwgC8EYOgeA9tBI+5Hb1advhevSo8g5Lw4AUNdRdxHCbHpi2l+foZze1nc4jQBZC2YqsXMSM
6IZl1f1hGN+9O2JGlW3A4vSgm6bEm+062AnsNJqeWKOhYR4V2tOC5EUVKqoBQPdMxJJJ846aphCO
PMwwgArwl003BzmGCHtmIapjtvv121aVl2gcT89WjJh29kO5rInjW912vVdpoVYC14jxqKYfxj7a
+FyBz9LSkuA0W6ydUzkDMA4Dzr2fABWalqTWVDHo+JxMxH26ULGJ5FWDWhkZHN7VYjJtVkUuOc0N
CY9RjTdlQIan0Yd7cehxoNvmj6ezD9Xc93B5TZxoV9wPljza0G3IUanbAcbIXvwsXC9hX5UD4r5J
N1VRWETkjasBPhZrV388cj4FZfUOi1ZpF4uA5YEA635HpSHx2wgVsTa0GFNoqGIGqnXjuQYzcE5J
OgnOzovTsQh7E8lj70n9JhR0dSEpuNeJDIUhAzVP8fkSZiVwwhetYWR8/hZKa2cqzetSXGMxPkDZ
DFZzLp2kk4odtaC3FAReEr3y3tagSf+kxhdg2U/DjA9/3bqn3NCvsekcQa/sE3Ke1lbNKwPAdD2X
+TGr5XyB7MYkOqx4uRDCFNZYPrzi2n/aXByn2GvkDBKJZA9q7NQCYbVjmaeMuHFGk6p1gRsPD/f7
NNe1ckjC9sE9UJhwCZTVFbTApij17pRwd5K1WRRe2INzsGRvNA3Bgi0pB+hNuGACPNsEuUnlT6oj
IBl94T2i7L64rjJDWhIPRVQMuoOZQtF1Cw2keBHyXaQpezl9loZBzgHSYYgXjVnkL3eNb67sBRfX
MGT33mZwR7gag7ZAJsq5/5sB5S2heNHQdZCFk/t8stBoSpiaUj1QDsDL1KbpN2HLoZ9n/IJotwOu
5KyQfjYlXLt01uOrH+m9Ks7T+209gOLBqzOVxyrg8BkZ31DJ7EnDUmshId/g6RI7k2jo8yEQ4lra
CuHys5ALFOxUKWM9W3RT4mXSW38ozHv5RtZE3pwDKqezXwepG62eEJGR8T9bcQxNiwaeuxL3WbhN
4A+FJH6s50KrJXH9CBTizpAAmyhrYwxnzAcBQC8IZB+0KmlqhIqfQZknXhG3mqwk2cfqabgmqCZX
2EDgai8c9AMYqIsKw8pAiG7fS5+GgXC821ejxhGs196vk+GseVx/g7awYNNNbSlSbYk1M+4e/75K
coQmlaue/AmFAm5XtamVSlKP5CglSQABMbY1w6E8KgaVixR/EW7UoF96thN9L5DnheNiVZhhmNqf
vRUPC14sKa2kziZlVcV1T2sPm+xJUz8kwcvDxW1B638Ou+Fm/j/WYxxM1Lw7XA75ILJdP7ZRcDst
Y0gffPA1kMhAIpRfPKBM/smYknLCBbyF/jiDzeFU6kJY2WaJ+yyQrzXFofpYkXnoeyWMQYrzEYWZ
0PCxM707f/rsnpZeRbFc2p1dGvb0MbEtoPejf98WedYLbpKd08myIdwMyRImuFwyuIIOGrgcVqTp
UMIJ/jV1ohOtFMkAUKIV0tgNRNSoNPcObN3yHkffbfsgx4pM/OEf9dIolTPMFF4jHfcpzl1R1lct
gp9GI517+y45HkwjnDqIFRBbwMTn7gQQ4K+FY+ahDB86eYG/Vi2On5/xX83Ew+FN0wZo49BvT+po
1+6z4PF8q4sJ3gQU0FKJWG15/m98kXWTACREzH/sJgLlwzw7+RofR6K+z8ss5xr5VNXu2yVntoTu
v363JuBIMgfgOSZRsyNQh7qmTqmzhtDMtCWtqAlRZS6JtCmXNmZIaoDG63a0evsiPhQd4H9w3LI1
rA25nVB5EPddxpiVQG7t81fiVvmaXk8v8ZnoAiD2BLA3a5bsPRWT4KXLM+OHaChfDgui9REkunxV
oawJl2sQegOhKEwl3D0RmLSUZvHijtal/K+N3DTi1nV+HqIH2L6Fjkjy2Mm1Ygq5GcqWj6imQAt3
eZkvECQLFDI715Avtgnnyhvz9r6lTZqneXPOHQG911wajdU/hBCq2C6CCssgiidxYSV5SbhfZlyc
VG92rJsnUxsphRxCADgEVCm7oP/0dgnnmSTwmZYPTpd7JX1iQ4+ZgD2i3TFXTjDoJyybPwqBuFQZ
PyHEqYlZnQydfU+9D/GmPpEDmkwhGkYGOVQ8xhja26dhL10myvDDhqX+w1zuT1F+g4SvgCgc11kA
78iNLM5DAOMnl7xjTzU1FejpFPvTIYWx1/Wml+TEdrjxYV+gRX8aexW+wTco2EM9b6JHNkOMHjJW
pWk6R0GjByo8onG0ons14WCJOFvlzLiOc+yarC14ixgbkEeC9JOGzgxrUpQzVgsCBjji3VLBmuHa
mi1v08Nfm44RCgDXmaObM9KmdwLaLSY+kytBe9+ojk/edZ9MP0sqbeyfkWdNuGYhjhwL2tWnXeyK
qNdL8NJ0EJfoi5N+IrZEqBkRAPwUTU8U2YmsQBH61iriMEf6iuX/lcev2ATwBWPH4XeFp/5CGZUG
NSYGFjp1mZ3DLVY+83ajrNGT/fzwQwmrC3NPcfgvmnmPm0w6ZRQ3h5lbjn27H86L7Ihfe9d9SnQp
T9+xHqoyvysS/zpVaz/5PzsutQFQ7H7uERVQw6oVvFsSnuacCPDagVLAOFK3JvRwH1dq/f/BGHl5
cUoDtja/wnC/u93m8VaLQjDZ9QFE4GCJZq9vdgIQsCNKR53kY0sgykGdlLd2z//Qei5s+u5aUcFq
BUymjrnHtFpDF71Sqmq3cUbuFRJoOHARXnWCJOasW6AOccnWwcyhO+ySANKpjAPXJrbwqhrA1Y8S
gUgVHGKFjVsMM024dnxkkkT6Q2cGxFKQCV3XNv7RFKFQzZpyl+fCVcRjg4dZFucJDUNPxlKHfVGE
NOrvGcf6mZRczFCKffYVkIbgUh/gTGTJRxuMFJB/LBjuti9NM4o9N0Qc0SX5R9oig46N4gpU/Yss
9+ulL5MVk70ws+cDhIvPrhKGO4JCSjNO1PxuPL7YXKhzCLTAlqts+mYDoa+m0Exjcr0PJ1P+RC9N
PjeW9uxjzDv4uPE64GV4979ptTLbEVy0QGXQS590ZMEFRbP1bbqv86EddiHeDyWQC/az9qBd6Lo7
eV+H/VVLvd16P0Lv+qzd++OSfob9dUoChsvQ7a71gtZzSIZpNZ7ne+N/OHiyDNL5WF9APjgxP20B
cRAIXQO4ijal4htGX1JHUOwU3WgpooCi/sIY4b/ttyxQZcwxxWenACSElWSQNpZVmMG33OhA/4Sv
9fzt5uJn57dfFYoijlnDVDFU7Em/Y8CmV5GhUOooY/CyIcXaeTZTEJ6/zVgK/ULp5Qdh45YeL6/x
JGCLY/2ktVy/mOtjAptF/0kaoYae7xGPeqhA2RS+5A68RVU23PIJ0m9ENc4kIpWvHTe4OM1hweC1
ETI4E8q8xrTYGi8NdY4ilyb9CehaKZJRlNw/B6cxOsVqk9qVaJO0zdzDxAlNjT78+kJYJTdnkJlR
+1pZzuo+SgJ6rJruOLOZ9ntoI+R4VEtl08VVBfeuRc3gyRTNk2CYv0nI8kH+xAXHoBh7JvXLhlHe
jGwPTuUfwSoLB+DcbJcvonykGln1uH4O6KpY36uaiINWSpEIwfDSZn5vI0N/ty0TiGVP08S4bbDQ
+G/ZUV+WLtTAOGYvlhsaDMv9X2ZqYrpj98tZBDLDcwnqVGdaFYRQin9JYuYsiR8JXj1WyqzBDWIs
BfAv4uWqqiu+QQCixrc2XuRjXq8zCwei9UUlMU/UcaiflKW8z/VsQQbvaNKm+g59xgBsiw+fyh6j
8A1EAahELpIxB3piELf66eiXQSldnv9mZ74DNndY9FSeVAp9OsFJTu99yWMDzevdLCMYYMfdvo6L
rsU59o24K7fosxi5q8F+i6tlbFRHJ6WfMF2KrQty1agngsJwQaDmTFw+mJV13tM+sc5qPth9mxn4
cf02p2g6R2plfaV3Mpb5HpRy+Cr9CHkwIRisoa23I4i2YusqspfLmQ3vAfVByB8cFa7yLEZTrShk
Ysyhd3Haz8a7VakdRULJsUVwODtGvUBU9WLOE28/Obq+nyhTnSQiD3g8i21s5kVJXiTsKnr4Oc8t
RBycjhz0M2Q+61QfFahIq85ALsVzDjRkR6mLO7XnCCK/nCzJ5CunZsXq4l86WOyVx76jLQViBLRm
stewSBYW3ltLgWpYlpVRWmHtQXgSZoKCekBTTKvAR0ThS/j13eymy8WxytKpLyovHravlr4mC22n
oNBiHFrOYPne0OYN257pNGmZ+qgltk8j2KwGlQW2ixzavJAdmjVtMBqEPhYKFKLT8qeautzrdtKB
9iCcm/C1hnb2ouxOOGA08rI2kSxp7w8vB5uBeqpqOwUJmu/PB4xW9KhaP5gTmpEJYnLQyN0EVrYt
R2SPMjYsrhaiU/gLqF2kCvb3JmmA9gkyAgaP6wWq4Xly7zDddELRjEhAOWosJ2ZXykrwQeEwpIw2
Kjk9nOAVaMv5zlFB66sVQ/a/qd5E3/OwKYyiGluMeR018VAhAZQ5943WzvmPgbXTZX6TGY3Ew9Jo
04Ld45m+Zk50lTpA/TY+jw9Oc2xfMheIyzQ7fcBVAAOAGUzLHJCdur29RAr8x/BOnhVqC7OZKsp5
pNPUIxqylIqPsN1buq1kAMYbOQ9bkuKlO4utsc55GjlHeI0fb+xhNjpLoG5uF3sSROve9jsaPsKH
1vXf2T5+xLtUQEekU2qHqyddySrZ0ZOrrfAj+xw0e2WfA7/cpARs9pcbRAr7a+wQEWrOyBlQ1Ngd
b7EYIij89/Te+upeGJCSRkb3tmcuxSoz+7kZrVf73JESVTZk9L1bCNnER6Gxp7SevImIR6M1aD78
H7lpm5smnDxNgMjs7R+eynBNNyszE1pMyY45xX/J0dVOcguBjUL1RnbOcw9EI3IhsQM2uuj0yK82
kM3ppSwzBG9pY52XvhgHtguq4SDelWGGPGRmt2GRceTZ4GGOTt0l0cXBvgFnGcq7+arhjri/GR+U
ar6/61VLAJFmEdmW08rtt8e2Jp1ersBsPaeziyOnOv8TsVRqw19nTc/gQ2z6BuTqcrDsEa3pHH0+
bTzQ8BVJ/43CB3XITjnLeg/5iHXBqzoSt72w8FE2Ewa0VuU0rlv8IFe6xptTJoz8e81g1vA/SGD1
7wxY+ZbRmcAAWe4y66PUFHWF8dUyXb9dsQYR0TA0pda5t2XxWSQhswolid2rernAA3PjoAIB2m5j
RlKEAU8klTbRZuhltyKqM9BHTuSG0uwLEDLowQHvjpmQXdDjRTvRhNcq3LyJNGRf+T0Y1R+J6k9l
OQF1ENWfsQjngA/RXIJlvqulSppwFcrFF/KnJhlst2K5hIMDegwIM/Hnnw9pYHcBUEAmgUMKNQas
qXjXQjdFEqobyFmNQtee1vnznFXBvMLvnQBnxbgauE3YZeyTdKaoQd8AgBlDzUdiCeXIEjhheBXC
S+AsaFjVKaSy3d/6GkJsW+evXr/v8+bPwudGaCWRkeVBXCpsxKTQ6cJC0om2yX9q4sJNODp55HqP
4xY4HANq4hcDsPXek4vUQ7E+gsGKkE+ebKQU5j3ADikzPmmS7Mjvgp3tgM0zFuA29/lgSar6DAjY
2NZkHB3DrwWVVL5FMTRaGjY3vKYaZwlzByvwPptkgrxloT9Ge+pomEFn5yQNmw3BwhfU0LpLB3Kx
sl2Xjd+HsQtEFVGlt6cmNA8u+Z//fZqze+S7llMkH2bgo4Q/Hk4xj6VO1fmdaB9+dMJprMkLf5gC
5ycosmsv7uTG1qYq2tUYBfBd1M2u58TB4j0dXV0SWAIJ3Hwyh2G1qO3/yV1r7ilppBo+bbu31d6e
JDnZByJ4brP/5/7Vzi1SjdTznSoozByxcfAXSgKYQTrNyO2PZDeMFMHJXrrLh1PmaszyMbLye/P7
8y9/6RoN0u1nU9/nUKb/wY2V5uWCMToiYG9+cSY7pnPwZSqIust5Mar8piSg9VVcOCo9JnPLvDeT
Sz3eUz4zhjNoR1MYk1rOfrtrjaIDxaHl0kNm2XUVnE02N/8cPr2+FkY9uKSs9pGjZtLXTvkhHVVM
ezfUA+wp+ZBPTtldOEk9eom0Z7hGy4526IMiaCMQ6aBagSXAu+mEBL/ZrVlvDmyBA6bhsinSr033
Z3pJfxaMZqmcODNEmAZG3IdkkpdpkcbhXu3a1coiLgkfHyc+dB0L87ZbpCMObnGH74ytbl9k7/j1
nEAvrpJ4vYLu2tgvRvXpufvi/VsYVwIsoybsjAWjdcUiBvnCP4v3ybeOQvPtqwthGxigKI5xGO13
O/fLRlR9aIkKiXn6GGosl8u/zP1JtTWosm1PInNLbWXU7AAOQ8v8O0w09EECpXCcGs3n9pNvksHT
/F70RTpqIWN3ojzPvtJN0FPWI3Lr6nUoc7VTw8weXlfmuNYhASZ/AFGF/3HU7XKedTmL8GcJ7gIg
UoZMNNnITnO8DKYQUR3Hfic637G8G54adj5Uz6ajHyQMGG/uwSvI/12meLe/me5SrlKRaqk/Ol8Q
Rw32agPJgzml8archt8OveVtbNwkjD8chxJOT/hKi6BumrPmJpjqOzzI1UJ/V/xLOvGzQoGbaKOl
zqE/gFsEvmPerkYppaZJ8eZImdcDIDVnr6/rauiF4mf0HVW6OMf4ieZcSFJqeKixxfW+9s97JXV+
dQja+QG05GaL9P/MQQeNVCsvcW2rhlO+9q0RlEExzS0ugPXs8Vc9hm3AV7+yZS+wk2pTDMfWPNnH
fSOGvywNAGnDrGEdTAv9Qgng7zv6W++Knhoh5uAPXrEZ8Snh4HoDSLf+BiU8E4Ou77USEdl2Kryx
dgd2txdOtcWN0xYzbeKNOdd5bEY9LGelAFOd15m6e7smjq+cpP0aAqrJ2dN1QDm9oOULT7/vMdab
zzgercmci/AJf+gqKF3rXZFZaS0ZsibNpo5jBP7ravS4RPM9L0bNSmbCjNFNPxGa9diwArLEGW+z
JaBh3QKMZwOnAQCkJ1xHfv/nvirMK0qkH0lvS8wsIvJ9lQObspgxpju7aQt/f5V/33a1suuTRmrY
1ANheto1iONsvNeyvYPWE6tnsZQ0a9u7uA+bze1DEhkwi7Q2jwtGwxiTgAbf/iaOBcMJwBS5wPiw
emn3N8OzLSRmR3ZscnCHKr6g8sW1cXD2DOIJi0T3pm6b0k78ICY4UFAreHGgU+CDmLfkVCLtL48C
Qaf594oGfMayCNAEnBXBkA/Tq1J4DRVTJhaxOCvgUtMCRFsNQ+ex8rZXz0GkeOBy/OlZuI7U6wWm
5MJUSt2WKBmapiytF1QD/RTCvCIL9XJPFYzP6wcwy0Y53NH3YuyKXMeYgJATqnokBvVtrbBAxEcr
9rutcAI57VWV7Z5sOLHVrEc2HI/MKeE8xCFZGiH0mtAWNtxTJWd/zyTwKq5Ljvu5eGoGl93nztJZ
0LVNYvA1AxJkXcndzPkvazMAWAAryG63ZGi5U4wJCUDj3Ygw96K8jkai0VmNp8SciUd3wjAE+2ob
q6ZnMCvK0hADRIV82SaLq9k3UDPLuSjbXCnoUyB98tUHlljZF2wc43doYUTAzy+AiDZdWdPxHk9O
QUDXhITXuqgb0BTRjkRnke/vWYCXLMyLFaoMIWN5IbH6Xg28qnvFkatFqXUQXMIyn8crHIIyX6Yn
75cXi5dTFJlvCOjQTqkpLXtCraAP4hbRwfiaD/VrORgWhOKUWCWLQBhNSzTC2Vtns7WLlXJyOayV
+8E/Vy7+ddIElZoivl1HSbrlr0PG7w9iM8bmzaQcNKgwtwLqWDbxFPfXwuDbAaf+EGfzVjl63Epk
WY4jcZSTxbId1pmnih1NinKmkUSSgr+mSabB+zJz+TduvpN5BHIoFoviLiegS5r3t12NdmrLmBwo
4ng0woG+IgI1KkO9r+5SFxt7soy7TtexbD7ZwEHGJ9M2hyEIVuIFOA2gfCJoHUbqg+zADup0EVsg
41izskBArLxKfaFGKiufjpbkwVt/9xegXcI9/s1cHi9OIrOaH3XVPdWi7LayxMr9iSATReKNZ9SN
ASxZnIfKVnyxGjgJ1rXJxQnGycVCfnnCntiFi5Ddea2pg4pbQrxWSqPczgM4yhlFvCDjS4W5MEZ4
cupdSlZpkF0hPmf/LpFpnoNLcRl9mNJtbj7+CrKOJ+8QAIsqh5gVGt8fuOCyzmLkPYS47o1c3IG5
+gMD5xaEpcr/Sr2ueWCAFbrmsRx4GmnoaxQnK+UlkEEmrw3F8It4sGMa1E1hY6zbiL7uorQZuGrj
mqp+VloUWGqVnsciLKbMxaiWLlgdEJ1g9ineSsdkWuOVOMWxDOKLdQaPaqap4u1BwwuXKyFnLUky
KTyif0JhgjA7QzY3NAZbZ79+JO8vH3D8XQeoXt3wtElH1fBfTB2B6U/tyfG2QVXBl/1wlE0N6hnI
ktBqQIcUj8KH14VHWY21v+rkudRt0LU8xRiNerkMW7FtILtk2s+Qb7x86SXXI7vd6PH/lqhtePkI
s/AnB/PJ75BRAM2lX47mJ41W1J0B5l4WM3oeetPxrvZLW18UpmjugoCPKDUAn73PFuaNZoGPPYCW
c3Pt4pyHDG545DpWs/l5pGTzSibSzl83K8nJd2smE8tbnCS/7b76Q9jDKevBekeH3aD7MANSGiRd
wTKpnpHl5xEXRW7ixNlxb/8w1iyUSLEaGmNDT88cmz3VTHzXSXPZ9FXwdJHljDGQu2oMAka9prHJ
8TiiHmAdfJrvSBAol+9DmRAmT3whoOkksNSq7Fi6bIgtsHc9AdQMGhVOILUUmFTfbDcdNP59fdYS
Qry4FNH49YJnhECyK3Nyt165tjKwcTwXKsb1F4srRKP6r4L+b9qqd7lURoE6H288BsYUvVR7fbDW
kqxJGjLyyP1D8UyNwnq6VqwQulvgrgp77gc/6IthZuuMFjdSzgi5wy26nG2e7vjj4WQuIhL9kxTF
IX7b9Ddcqwdl26SjAk+aqTe413fOUoRsakZ6qhNy8ByIZQrvSPhGh9gVy/1CPCtLlmxF6qOkYBOs
pYcapptospxAgF5vDVkwNkLpM6GUV9ggVOGxPsae8J1LX6JBVqr2beDeZMS+IHgaPZiAiVnY91qG
kK9lc09fkaCz9RbbPJlB2J3RqadcTQczNmE2rUMuscYw6TRKGsacu5gf1JDAWPk6VR4y49YTjQ69
EZO3fnfaLdx4JibQJBhQlVM131iUi6ncfNCUiB2D5FTIuMcxhc8O+K7PZn9+cSlvgeWzyNQaVzca
QVVxw9CkJQazDkNP0knkfCClGqOA76m+xyK8uDjbxl56x1gTK/CwrVWHWn0GFM7knFzZS0UxcrPL
ebYoH8XyYmenkF+xDp7pb2kadDKzIikwau33H0TPKjGjS623/ZvRne3GNq8p9j5UE9G3shNzykD4
K4EuV6TmwT+mfgunudSOXT65okyHZrPQYChiv2h0VlG/J4Sc/QWpQ/puUztkEzYN0MB+WoJHlBiF
U+7TUl3nTc3KI2/xNYT+c9SIgQnEEANX6Ui4mNaeGUFFufYZAoPupqlr9K0hc53StXWAyzj5Blhy
ib69L8cz69EIlDvPzEZY/uUL31rmf0HbwpBhgCN+8HvNKrZ6Lasw+EzjxZpB+Je/dSCZ2k4UtqcK
5E0tvm7iWmwuKOBN91S1OvCBuJ5JgsN8gQKxn+GzaAnMM8lmvBDutT7OVsGQy4k8xAYLYb7K2XTD
KFKnNFtKWcFxHBGbXOeuLf1A09vRQOJYR2SM1j0NglpFqTtUffQPNqCa/FpCBH00C2xgoVcYwFr4
9KODe0IUlKFUepH+8Fzwan3WBCivc17KcdcqbXk8nJIUa+nSMdBt7FznDycAg+FNXCmF/AFMQ6jW
P4il1csFxhuhok6+w8kwrSp2azMEpzc0bNvuXME1PVHbqy3vrVZE1sctUXwQhMYgPBJtvmVKc3M/
kRHnl8w2otjiXPZPnzQrAvrc4TBMk6jfUVKKBdj/u68y4ZYcQ5SgBGvsY7Mtis0sqe4EQfGQiGGs
klDew8xsJJrjUqGY1P/zJ4L9Sv3ELQJMQe5Cr8WIay/POuNYmPgl4+DI1ftDGB54VEvrm6jJypP/
MePD/WqmxVRyoscuSCknBAFE7qhSYMCUotBSE2dMWilpz1JNN+Of+iWjJCPpN0PEWLiAKjHR1g17
xFsMAoPb5Q9pWLngw5fngn0zrfmW2JKaojkuzBBaM3axgaLgzcoHE4aW8DKmSq2btIkrRqux+NBJ
of51nRI2OxmRd5dN90wu/jNtce4Lm7wAo+j/hTzc/qCeueKGkgYb39CfyivEVOOukZAdyZ+SROps
nWDBga9lT6geBClCgscT6I5G2XQBNKw0hnsO/qJdkjSqLMM0KMhVIV2qomOOZ7YVixS61phKLMox
/wxc0WC8tc0qHDYXqnrQgVNBCEF/IetCgDMBk2kvSPcqrS5ipFO5y7bYzMq7K3+V+yAetIAbk31B
lt3TSEjxOlCIC/qSEKU/sK+gvLMzz5n2aslKIgB/taLcQMDgR97H25iKXy3mRqLZCht8PVa0QyHu
Sh8HqRuJ2Xy0NvWUzI1c/jUlr8peAqlIFoi0dYu4JbfpAuohXCvT81GJmW6D1lpOzd0/mpwPzP8r
jw69Yd9IKZJ6UpF5uNLnQvFbnIkqVkIWBX/8nGMW8TiWx0rNokyM8ymjlHhApyFaH5zL8w5UNYe7
BW+tTVIVQr4NJFEUKwoRdx82W1TAVaMzxmpnJw/TO7vYksSv0jjiSbd7tcU0J3XM1Jyy/PFHQpOp
gW/Er7dfkAeehHYpqYOZNfUeGAyxhjnGAF0xAMpjViHHpnpMzSyzAJ/oQ+sfoFNP3GSMcSgsCe0t
Xe5xjD+ZR3dI4R/UlND8UdnSQK21ZhmcpcKGC9vulh/J6gaP8I70fua1kQF9Z0C6ffG1vK6WhLdL
nNrgJAPJ8V4jdsO3TbqZZKqAtflgFyD1O5EKaoTAu9zslTPseeIx/oNA+kH2D0pMJrpMc3+22ejV
b/NFGXSLy7hdgwqG7vajIwhTHql1K6Uz3KwcNxzzQ5u7Kq1sJ5+LhetGhDhEBQDix178XZMwyXqr
e/joD1VuwKKEy38vqhHYS1ZtAPFTHXGcCAUeDB2s+6MgSfOg2d1ZP6cITQgMapSp50/1703OXGcP
UuC82aZbw/4DAV+KHVJlg0QEVljZmLAEzsjaOdHd/vF4Bhk4dgfPsRvyKnjPI629jljWOZ5Tz2kw
pFup3GvrvKojiH5eLf0ERZc8xcjqVUBOBI1JBWSSrqEWuvHY7u306QctZwXEqslvY641t6K36bEC
fzKTwaTrMh/M52RfTr3xVrbaafcPKc0pCwOZ3esW3bkLL+219RywWfOd93SXWB/DmsKDvw07s07k
wIP4wH57iT/gmVBosR1DNIQKNjyqfVWNYUCQ4GQfNSol40d26EqKFpDhtlMjdcq4+P05r7RqGZZ1
FcOb+0eYynW8udeiJ53AA2eHCR3L5hqfn9AD9ukax2gpV3Z31hktQSEqHAsgSKCINkJ5C/ANKvFt
DtLdBJb8MoFbUYNdlyl8C4D7+H+6sJP79wWP4Vbm0fNG/tmia+RXgkbVvZg/dNhzzzhDBefhBq/k
ONkQlLvyhLc98ylhRF6Ccm62wegnJUyl1J7E0J8pWZMphhHrY+L5HNuUHscw9ws1UnDN046lYnRx
dvzgsAlWvmya6yL0cGX/Evdd0hFEug3XrtzWjdXLZPHsgyhC/Qi7xlzOrVMLsWBr8P447lhuqp9w
VQBmRAST9F14pXD+dKjhQFUbj3glmCkmfpk5casMhKM9C08IPFmQdCgdyFkKjKlOsVs7ZJ3k5ajp
+tKTbjbwU8tQnPn7wXVcw5Nw6Vdx/wZpaFrnw/XUHECykLMo/vhJzogwET7DiKiNacwvDv2wOAeU
AuEzMEoMlHvauKDgrCJL1AgnJiUP3i1eEUKJdNIhOAtym+O2hH1FT/5Co8kuf9rJ5FybO4Ye8tg1
w01t4A1xgEzrDlMEREJ7FOgea4ZzGjh5M7BESRww4iFzVH3LGJRD5V5JL1sfp6T9vfIzO73yi3hH
Ze+ayEcpYsINeNrUfCVfdR4LhdWPVd0tP6gM8LkIVEHb81cp9ZYIId2+iJSpw/VaddzdfRauNNpd
ntog7U5DrWfPXTBCibo0fzuqVLXZ1ghePruyE5XaPBZoTsdti4+ed2TeIpPxx9fC2rR4UG6lWsnq
r7H0gO41qrnnDIKC7iFiCl70r3XCJEeFJn1PRQG/hdDDBUKjAoeQa6ToOqAsIJ1FmS4x4fvoKdqh
3hIOfUT77Z0caQc8BnL+TFh/7SygAXnUY0zZErzglS6lr0MoYUrI+7poORDs6e8acgsmukU0NhM/
rIKAxY2tVtz25Htd383cpmOYkvbOMFDEzca8W8ndlC/qa2UGWEIFIY9aw4yus8bVdoFcs2Lcbe0D
09Kn8wWyJ7ZQ+Tqr9wlhQ/QqAhyPSwSCcnE2S0MnbB7K0GQoR49rabcO+4zAMYbEaeve3Zn1OjwT
r0mdtsy6fYZGJ7kuhYI34G/FP/xvfYNKE9ptRNNEAszxi+B+y2fKZFL5etH4wo0LXlyKmITFimw1
/BQeMQHv2zgL5TPsbaIEJWiMY+U8/clrAdTYjkVUWWrddm5z3mncfWWD5D1NgZtar9RfmoJjGIgg
qla5+AtQmMcwLTLEoxijFAUQ3Q+GVEE3XO6IkRvQhc51oXo/vp483byV/xHkLCK0XFGmD0eCaSyy
CdolF5QMToNEvw0fLmw4quVFuVzM6rVg6TtJNWaLS/vrTjNhi/J+SGDc95j7EgaoFYBJ6St5t2li
huZWy0MM67aYWk+0by8aTisLGxKVeiDxhv2NGo5bHmaAl5mHM3YgptEUZyNXSiGVrOrr2DZPJ1md
DChiSdQ5KD492TstaA58udWc/YfbNHKrNrUFKZHIOCeaELFMtQFX9k3SlXmq5Ztz0sNurcL+Usqm
vsY4aYBZJYm47bjI6K2eobnCnGPJgtdlsm7ZHbbPmXqkfmL9IBTThVywwDzV3g7MksxgZCv8aDQ5
t6NSq3+kXxIjqutoIebwtXBJB3aHk4luFSmS/03+SuIGhlFsL/WuJPwWXULw3mmtqtWtFKTFj2WY
LnEXYDTFcy/8vUs+mI+pg2ScYKl841xWAPZ6ZQfODK5ADs7CdRS7NTDrQ2xrDn8+o6N+11IsFsHO
QIZYGDJECMzwG5Rj+gIiLske9K0H5e5DEcuJ0adQshDLMawAeMQNDe/56UCKlYwaS5HcNLDWsReD
tEHrPP7gBt+di64BfGMIE4seiE3khblkOIN0YSR5LdBAx0uSO7E74rXvVExgjEGrNyLyMu489uBp
eYX5t3MsQdtZc0xjHYoDpmsixa6j9sPZvGRrk1SuSLHFjJq8rVUF7jTDixc2PzzyQR921J+uCWX7
fqyrRH4T5J1S49c/Z/NWJbl+h95Te2XSJo7XsFK0K5JTATkEYMEShBFKS4mfo8uKjbok+IIle4hF
LRy2Sa/JCwmLWlf8VLCAyoQoSoKulnqdfqZB8AJfu9Pe9hCY1Tw7/6w8qhMtznitBs3Em9VvXWPb
R7pJzLEElyFNSsS9rLx36ZnTChYW99Xou3UBU+XfZrI4LN9ljg99K/zHp9t76sYN8O0Vln+XjrAQ
mc2OV9wh2IIUPbxMuZwyzXENvq+JojhKHp7n4VwY0xnrmZ2oD1rBepfkjDkS/Di2YM8nBa4i9jG1
KJdh067y0y3AQ42qKO6Qe0ESWf4GGAzbvnUBBg5tKFLcjLc7YneRmH2wdPF3l/Yt0WI6NunaskEz
f703h3BFyIz4EQh4Jp56OniIE0rFH8sLcQFy/hj9yP/MwJQJOmQds0lN7j9LhXZ4TzSIb1y8e/+9
D8Oe1jXtF+ma6MmmePagZRuIx0ke5iLWxGJEgcVn4tWhYLTLmew5w/SxIs0vSKEPlyMiXWoIaXJA
EZsB4eugu9p6PFeRU4my5HvzF8dilweukm2KRU6vYp14QQfMLOtNJoqMhvJ+DwmtDcsh7vaP7GH2
P162Ue+PLsiKIDTx3t2spN7PgjN8wXscAHxPEbVp4yQadYvjeXE0SzGJiAqTjFN/unl2PPixAU/z
fWA69onsw70SC/OTpxSlTtMyeop4MelspyuUziArSVXg5q2FgEfQtUBha4CnClkoNHPJG+WpPZVk
T6YHYFyckfZe9DsyS3opzux/92knRy9IKMhqpJ0RVpcNxpkcCyXk6O3j9wuRrzEFouogxyvwICCr
GBBheDwowmiYtuwjqUCq4k+/6iZ7F8aOLK4vShSxt7OsBld0XJPFeoZ24tHu1rZ/dJETGx2mfB9I
yp/2HajUi5cpGsRXoB8cNlkbWKCtSApIAlUVEZmKEAXfEHgM/KRq77sesK41nkChcXkm6Xc06jTE
iiyw+P0Gna/xAP5EcQSnxXT7VXLFd3yxUnVeTF9zlRjEX5iaSfs6ZITZnxeD8lDexhAH1+0rM+Kr
h1xIKcNdRjDwGDTXrnI/gx0fF6d86GiXq05ghRAdn7Xg5GtodVEJslzbnv4oKHd5/T6PKpAkg9EB
2XEjnuj0b4UZmOqvlV5RYvidOCs05k1FYrqdkA9jrKPtkCrfPBrz7rymScOyFIf4L6KJN/R6I79Y
ECpkTj3yErsmA88zGWUjZCx3ybsNnMmYlOQcaTBDngKx1oRt/6NQk+NtX+yQdi6fg9HLo08CCem3
oHk1F9VTMJYQw5FKhAiUrMaLw8Vst5N57fVu/nIq+2sJLhdzBqZD6Wr/RE9SN6e/aAa9LeemuFh2
/FuVq7Rx8EiPLbhrjq9BTbIAIkfxMPaRNxo/QeQ6A+P68QXWzUW97fFJShKhS5LbetRpVLTaaHtn
GisMEUFDfOT7Sux9UAI5IcKm/EmH0k1vlU+LC4MKqccIsV6akCtEXozhDlKBoT/cAo5yJ/Sl+vIr
X63mU3IiCeCTkIlnXSzpW1qqwWsPcsHjrNU33xVOfUS5+9rF0ZmW3fMhUqP7sYi2iq0U1us+zsp6
OGE5IWjjnY1eZ8ohzJkS2R9bG7jgiKWQ8XfBwubLNAS6YNNfTyqdzP7onFvNBKqOHFPnStrj+vgf
1asnKnX+DTYf73odtW7gZklR1tSdT9a7XMyrG0Lz7rWjQKIXCWkt4fhHmS14PvM2IAWZElCvG9fd
7FBNt1RAg+IP342YRVoMiAEAQO6DvY2VQ8nnorOqDw3BG6NkkZAkl1g4Skv3uzXwxZf8JoG6PHqD
L86dPMen00nsc08oOYWxxYjDXbhcPrfPe7wveXIdyj8eBWU+6FdnWpx4cErHIOk1u4u5cZXXCz/0
GZFZvTTsBNpV2PvdNSp4fRqWMhqud9PCUnAxBqvbmKMQTgymEg6dTNpqC2adUSeH9Q+q2Xnadttx
x6t2UK+VA1Xl5izkmeNEG7XU7I33hEx023JCpzi6Iv37Ok4gKxbK3isAe8l82qmcUgBNxCv+iT+8
pSI0wIXR6WHJsCUETFAyQ83gKkaoon9i1uiuBu8YyE9HCrmkY69XnkGz3mtlIJtMZvG4DU+y6o4N
P5Qc3v8+5x40tp0NJI1qX8r1ZbKfsOZucv1T/wn8o6fywcKBJE8+T+POFm8B+KiJyqcclu410RnP
Q8BAi7D7oIVGWET3udXvS4CfE+PRkhZ231nr3FzMuREwzye2PLY9IhkiAXjEco4hQBhqAd4Srj8w
O6HTjxJ5N788ui4wNOkK+jOCCr4m47Utjd/hr5i1JaUquI5Gp+MvggYkLXYCAHTgeGOX46CmaeLt
otEEDJjJhVnoFCxLRTMxdr8WuQT/S2dbNsP1G8ViIKLu5cV4vGy0cGepp7UTpFq0RkonftQ55eeE
IJNkd8F984jk/lxWeVYB+tQsrU5SqoANjXTL2RFCKWUdv8S/0JY64x+P0h/r8EzfFKgvslucf+hB
KFoq8iNdWux86SScY1GMSZ5/lPWaDk8V227S95jlmVT5L3NrvMpbCMbiJmsdcHISoxBxk3P51CGD
RJJkTaJlt27dYvb1rIW0SFKaZdeP5wVh9oFg5YJX9lRwRXzK3m2Ou2zO9gSID1xSPzHUe+HpXhdc
DRsy78Lv4qJINDteuL0ZwnGBtN/rlyM+xqX8sADsNQIe4AzqvUpFRNNE9J3QnSVxrtBlK3laeVad
pTqGo7AaU9OfiC5MXQH/kNIqQw2QFGQb4B6rmO6bQNYs6Y6excMKbNagpG1mcp7gIK9qCdhvaJLC
Bhi31jnNrSdsEFeKGyxITrwcRT8PJFLql4VKF0M1vHKntZ10bFal6CFSrEhysrQyaPpLmmFae7Ke
tzC0I0epoEid4UcW/XAoX7U/kZnxq8hlRa38Y8JKDmnj9ez8b7kkV9ubTX8fbtOnabm98YlWwrHA
zVObKnqoHNwb6oe8iSjfLfFRRChr1Htzk8NT7Jd80V0J7lm89ATy/OF0JwfJtIYMoNce8lzhI5s9
0loYduAxCEBfiYeyJs8on9QMbkJyHYq7i7Aw7K6+OXZyX0Cbu2ujnaeH+l3NyjXbeOOeh8YbHctg
nhqPS82A+uwtNzywO0M5Wf7WEWAZtd+bF7l9EYuV4TOvPYTBQ8V8Gn/dpSBE0l9oqJBi9aKDuRze
3CPurhywU1aq86p4XmWdkTjcn7froo1Ev5hloB1Y08syqzOhvZ99RWhBruj45zDWggFLjrY5/jWZ
8VIfCocimkFeVhnUJU/0xPefNIG+Mn4gx4v72jNS6l3hvJML5TV0jm/wTHSecdbaZo2WmQNPqbJt
R8dwZN6h7MMRIgN4zMNtifbaANmF93wZa3CdMSvZGtBIK/Ozsag2ATWxe4uSTnC3dvfbe/N+v9fD
SL6N0dSiCfstX4l6l11hHHMubCGukfEpCoO/8GQxjn+NMpXXzHkMfoQ31Gk7dZ1MCf0erTYJsC05
OAd1oGTrYc/Ok85udoyvs4xWN6g3VVDwRfpNHLHjwtxYVSeuYuoR55x0B65A6u9dGBV4ctdlHP5i
+Dzxvwyqiba/63xSsaxQm4x+/MzeXdwKBx3IgcWTKFAuvGoJ5aYWOrkcuMWNxN7mdjl3Q/vq+6jp
w8ntE6S58V5rvzELBLlpMrR/dzZFcay5N66JBWQHW5RONO19KrQCtkctiHmMoNSvmE8koc4kLP9D
ztMHAdxJ9NZriRhYywaUQBBibgeyC38koZdkipOHkjn+cttM9QWogXdNFtynAxKGOYufpJsqvoqI
ZlsoVA+qZpoHkxCF2lCYqpu8j5+BocFblFoix8t0ArGCBkx5sPMscMO4N9zJfbZ1SXwbSNfgTbJd
gmaY9l/IwuflqlcU+hh7UiWdafEdRsYR1G1ARjYA15kJ6D36ieGQMBxPcn1sRxwdQtOLAhi24o0Z
9Tui5GsZqvwOmU7eteeEfN48HwaNoRiHaHEQC5ss0w3B6zLmPAfvUWtPiJkbYD9LKBX2fkumwCYJ
rFY31xkp3NLPCPzAESAOL7j/gqNqQkT6vWrYBOilR5cG/0DIouqglaT/xmHg7EpS0XOfF7UKA2tm
IK3QwJ2X0afgRLxYbHTEcMq94A15ZoNE+XUemx3Ro2eRqZQCrNiZ2mUNRYKTxISITGcRkS8RmfU6
jozXqroIbbGohDdyYffag780l61ZW8TbNBrI4PKOIQqxeH6qJIpVAKnjvo7iI0FlQyCp89iWQOH7
2La9lbp9/s0F4/mZYo0qFeT0LnSKKP1rXCnqXHH8A2V5QnUeQAulhmnMPwH+pebj+a24KLzd7ma1
6Wxk2/2Z20+d58uDmUiBMSRWSU5tbA2vPjFeFTEkpIFIqBSxf0vPl3dev+QFIUbCRoPpock7TH6w
TXDYqMAOPsc2ADAp3+lOkv0jOR61zDYf+WyEt4w3X2+i5rnJoIw0dgRBRcfjzePRXLmdhwL2vdGZ
jEjsT07NCyugK1BXPk0hhTW7Fw7ST+HoSU4WcNmthfZTir3xbe5iY3ZZ9pCvigb665Ey8FO5KKXG
+hKN9m8G/z+IMzX/vvZ+nkjss62jqcp0sbiXeI568aCYvMOD0x9raLZ1xpfXb/N4KUWN/GPFILKB
1u0Aq/IiYzsXzMeKgqJbxHPsJWS0b+TEIxYvzaBMQMDtBHGzfZDQY00I7Qki9HtrPsT6K9cFcgq9
bUugLGEzkVUjtZkokuP0X/DgO4yFlMHOvoavpE3qo1d5J2ROrNjuguRUNzcWDRQ08qhj2t12TORa
jRNoXw4TmC7+HCySw1K+l+PhtHwP+q19l3AEcLeEsjmIikjX4/yL3uf1dmyrpCbPX5qNEDQcDpuN
tpA1nGzU7lBqesjoGDHjKdCZJvIQZkPYxnNUmY42Jd3m2XtHpRZ9yJHDkMAAM2+NHm/vLpYqfHzg
rY2UJQvgVHl6zze7JDaGYAdqZjkyqLkbMRq2npMlfVJFG0aoGbGf6mrDoLYm1rqeBQQ9qSWzcqr4
GdomAsA/LCq+EVRHvGqIfvL4XcsDUzYludCc3br/okNqO+RveTdUkpSdCreOJb7DbZnfMX8h4h3O
goqUJl85l7lVDa1xtGLyY6i/pAtiei2OwSJzuJKyHE9JEZ9uGFqZEYGDy20qKp84bQ2Hjiuih0ne
myZACKkckEPRGwEFIh1lGAzdhfiAAqltcwqk78x5eLzgC3K8dlXgyz5utTV3SRlzYzlbWG7sUKQo
0g0A5v8T2oq/yggGfOYo9cuHW9O0c0ZZJwRd7MlPkoGKC5sc6O8xMXnnfEf5hF/9knskWvYdJyMQ
5PSdPf/r0p3W/zYZOR4JWqwst/vKF8o33gJH2veumSUTJIeS1qNpopOuZ7Tlrxbi2buE7fR93atd
Qths7YaP5G6WFR+b+mCYNBeKvfM9yMjhvk17r5COVkEi3uD9W8jeLDST9z/m9coNYc8Z+nrP/Sr5
kE5cLUow7MDd0XQvQTEgvHLZ9yiJ6LHx6t1Vud7LXvavuDRp6GbwP6JK++VcU1/Q0mLNAr6um5FV
QOwCs38ZAP5EKc0dOE9dW2iVP3PVPzjS0cGwDKL7tn22/uTP2TckaMm/qSNrAS7Hor8DxDIEI7Az
b/H0Aw5h0b4Wlhq6ZAFlG4hATrW05XSxo0Ms2GFexWc7mMJna01e+DNgihON9yp4V4BBoOt9wHXs
utMgKWeAFdkItnTmceMtM0OlNlASch2fHtp5Dp4TDz2GJOOGIk55v6Tmf/vXX/TmGUA6x6Ss9kIL
urH3BeAaYE9fNqtgH3+Jl9EDERle/IIKPm3SKE3VFVj/WUybO55Y1NcEXwUbYCLWPwOX+2cVyOo4
EhFQXXiTNrvB9H74eSt6WxO2UfC0kJW+xO+ihBq5QL+tWNzF9zBll381jAuYBv0W6/NkSpDfjZj3
2hyuZ4zrd+CVl9eqQ9OsUZEDyjnDZPdcPa0Z00fr0bijc5bhf5zoDTweOxMVHRrNPS/iLMkLmQvL
us28fLLPA8coXUchjZqehOd6jroFRbcLozI5qDGZJtiY/5D9LtBvVqttTPj6dGl9MEMCUhP9mfvX
WJ7vxkZDm/0NjggrPW9KWkT/9fk+klgUlnPvEDhRA3BIC64BlRv1Z7IKJLLQsk7eVUxi4UsRMi21
hl/PoM2qbdhVzJbYd0w93FUFbhRGQVX60dbXM8MX3q+VWvF0F6J80LkdS0V8q9Kn7FTSyZwJZZeo
ZmBfBarVYkiy3tGsGUqRqTpARJo9f7HAmnOF8IaCqz6abh1VnvnoLqMbwT6yvbA1EUCl+x10nn+u
fJhBnZIIYT+l7qygks6AOXiG1HDfnlsMsfNOO0U0i95nezqR+biFozgt28iXmcb9gIScXZAb7AdF
xlYzPwlRbtDLfz63edePODB07sqa5Glz4qecrBSCNjd5Tx0k8QO0QslrFjeT/NLmQ5mGiqLh+iut
gAoJAo920ybA/CqWX1K5EpjV0gYV+7xeWsg5oCp4vS8izilzlffugzDc3E2blrnmkT9pW73rbG5A
eIHfwAidL8+PINU9fUs9zHRpZ7mVbvdSUUSttSkRCejpJw/6GU2nkIlXSfkIddgZ18/Vrgso9no9
kUmZwSHxKcI+nDNXnJPjxGDTFtSyc7nsS04MNDtaZDKsYycMOP5F2Ot4ewoSIYVK8I9TzKRE5VPY
YfY8tH0ir2nZZPehyGN19qtJx2UWF4UGfL0sSw5VPVuyYHCvr+n29wgK49r69i5+z8h3Xmy4Nvxl
I7FB5ywz5wdPQjD6tUmidjnadu2qR3lGGOhfv6IFZNyAeY3LWy+RT+oS4S4tvhZPujg9J1YMiKNQ
U0cLCrYCyXX8ZxoP5bmYWPNBpB/W/cFMak4h9W4CC/ACH+qujWcY3CRnnd1j82xXGhuoURz9NHYj
ff4q8gNylW4cp+wD3rkXTLp+f4BEFeDFKrzhn7Wto6i/j2hk2sx+wjJZZcEEjIGF5HVxhdpmNsA3
NiA4PJtdj2OqX0hgBLlKJnhPKnj+3BZZ1DTa0xKuEceywTt39SOUuwFuBui1K/TMMAL2fSp/fTAy
NnRD8lCGT74bsKdUP6zhyvgKtYwi87eDiHwvFsgy2AKmUcX2k06QlqS6+mBgPc/I9CpzMYGJZiEz
O+ktLsnouKcnE0XBKR2u/XcQKVkr+tp5BXdTpCAWH54Yf+cS5TGhH5i/uVYOcAELUkFL/p7g+YU7
niUvmX+hOzSHzYDTQdJZYcVX3dSdHFVlU1B9pIuzYsA4y5mMv4nY3ez4JoVKOK6fQYS5Sj+jEvVg
O4lAGcGUrOLYrQw8nHVWeTNX5u8D3M9rdOisxZAG7Y6vsIjhwCix7hRye9vJsnbi09VDMHG41h3/
ajuU5RmfIHZKaXUyBKB4SDGazJZZlNJ0o09JVKzq7JET8VcAO0WOX/Bz9ACi+atDTBAaXPSrC9gS
IvkygdPYkfqQZBOt55ZFBlNp9avmiQeLTmsjK3F2wMgi7WPvGgtmm7DVxt9/5XjyoRjWAZGx7iCD
vPqBCIhCudOEI2hQajaBANyVsSoQ5mvbaDUZgfaPDTMP0csIPECW/u/ah6cisUtis/4uc1JvxAUD
GyB/dkOO1CiIH9bG7brjnED/7GY4Gv+fp+JmI6fqjkdotanjqQX7bUQDY9ggelLmrfd9TMS4NgdR
OdO7V9bEHM++wOpAnqUJxLS397O4s82yDSRqWO9fmlSeugyFHXHM0Kg2S/yj+52aAvCaon8601cC
txmAc3mKDS/LVvSYb5GMfkgx35+dN+pWfHS9qChWq9spOPFE/XpDOIizfXm3HCmq/ybyeyw18shr
SpM+XEscM1U7wVHcOlKgZzmKHnX/+x6l89n/vnAYGiJvqQzc+637DIbHyhv0AJkucdciJWNF3sAh
/7r99vCyVPdUQjNYYpx04uteGYnigfrZVa2j18Fyu90SnFveroWw4amJPJbUdrKMwNvFu5kwDUbV
VtmHB2SOnwsKtcGFbbiyR4iDO/aeb+aVxgSif/ddjGALUzjipbtDw1fZ6kCOr2OKo7+CF7eL15jy
z3CTuFfhogP0Nadhz1FVSuoJEovzPCSFjcjPXmLloLngyKuv0H9xwUl1Fr80DV5Qj8w+I/tO+oSN
l3A2h80suidLYHDfn3y69Cdh3kxkZFwe+CwbPRanEQdE+UDi1TtLghIFRFb9c/Jw5rY2U/JHQo1n
5TQU9ebreQNdZkFtZ7Q4iBWo8GpXsgwZLQZx9X5QKFS6Z093e95k2nBKtEP3gHPnrrZg7pqVDYlD
ynowt168VqYfDJqd98uoHiGDkXeq+8Iz7c3DGDNyJkqOAtJxF/tIzjeYJStYhjyACqCjLjYMfCkd
keG0Sb+IU3jUpCZ6DOhiOTPtIny8H5RVeH1gQ/shEJvVdjm37MDHZiCdvG7lEC3qZAGs2p1SpNwI
JhNXY8zVx2fK2S8VGKqB6SuHRt+QDATVlDlswAGN7tn8GfGivXnOavEAwJL41jxam5XBP+v5bLZJ
pRjun2fdLpOroMgtNrLVD9s9FUYZ2x8who6pRdB170OhfxdIT/uyuAjMumAs9mMCExbJuj+0v/a/
fi4Baln2HxAD6ZxFb33Qr+IaIiA0B9E+l2QMN4h4Iw/GCYyPRBKYApXevtNTIx1upK6fbIVYIM30
9I65xGt1ZRr+E8Szo/Oa8yyQzXFObBgRPsgT4Qz32sFhJ4jlRmtXYsFZ1dZVHgwm/SyOl/UfJW9/
nLtb/6CLxSqsnC3EFqvjs1aB8DqEN5nU1iu982ky/wL/8ZOGoA6VlUUwXdy+8kimrruD4xNA82er
bleunHWxqg5UriG/peeWpVunddlkriQ6YcN6ZmvoDYeszNynKJzmDwnFnU5IcFkk5dyHikC1/Adx
gYjLIn34ntIKhN+RPSazPI1rDRKdLowgmZK5ltmTs3MVI59qpOmRPDGNo0v601E909bMcvRARDcA
f0K0LdW80PYBfd1R9q1xkEGA6Vg9AhxkNe9iYCDhx60sEMmDdFU7KbFpT+IoNNPVGOBLALhA/TVr
A+XwZIYIoUJJsZOraLV9tYtcj1flWjfqnGM4gnZ5+5+u26cDahvGIy+LJ8h2Jgx2DCYo6F+2zJVR
slm1SrHWUI1ueyb2cTwZ6mm8hTmvxTkkFVWCW5U9h2d+iS6xVXs0tPjsLsufpunf+vHLElWxa9nj
e7PtX5T/z+dmdZb+y0mhBPgo4ue7nNBimhYxpzuNvR/esN6N6BNw0zohwA+Jm2dOCdSR8phbij6y
znpTDQbS5pwXvvjP2AatewsT4QkruMqxjIGgjR5d3ZeVdxgxeaI5fUHU4UD2oaKI+H3x14N6jfDC
GvhhjcWBjCwn68+YB7ImanFUjCc8Wu/3bfOUgqOS080BWN8WNgjVzKj+WJeMdD8rNmGLNX2CdGQ9
towLhr2yw8gQ5+WnqWVs1eXnXWm65x3ISX7PU30Tid2WNRsIDBEhTZvIeUFXW4UZzQ/WSzMmlJWC
+TtdU/IQTQdgKQtOfVp6nvWhGhj0auCIS5J/cXp84StoTsiDo+b2ACBwynGErbAmMjh1863/x8il
F1qSoJZ8XUghXdcll8TgJ3/XXMCVxT2/x5/B1bruDDWzyEip3HKgoNSc22b3uuWt3v9NN2K+jLSN
x14UsEb6NBgbbO1wgxS/x+eNFyXsdzqBcjdF6COmVFrU/7NEDnTmRBF1PU4X3OzztMfJjYJCl53U
fbsTldZsBV3SwqD7krlUlUoOhcQRIvEx2IEYYvE5heQ9UAVyT0sPDXTtvE/R9OqydzSvRcwyaMBN
R1OmTjea0G8FJlt+zTC45zL4O+kjyfMe42yB42YGs5CinF7jjkYsGc8ZoHC87QgPAXt70ZGjUxCw
aIaR6VxYn2X9gseY8B8m3RAnzv7w88RTmegUUJD9/6I1e19FXlsMb/E97sBMCQg07jO5fHJhB/CO
tU7EU859sbR7v3nrZWUh0YsnmiUVuh5XdzVhHioeTF636PkYjQugCoEy+57jmkFM7oW68vlnewaR
GzIOwC6OnxCSki+C0lbp49xGsIa9z9tFYgd8z29HZK9YCoSnb6fe1UJFIrhpfjeUwd2NLFVFfWgO
8Ys6/+HjLsL3i57mo5mpuepFRa3npoG7l1wE9VkqEfUTjTDWK9EFlG/E7Bb0R8NEB7U1Xdv022lZ
JTI0I/BT1bR73Bg890qpLcypOzxfO9lIQmCvPY0D+xizZLAv+DDJ5pIZl++ctoT62gDPZtebtuX3
EMIZ0E4CgNX6qqIyb5jZ6v1BCLhWYr2k+Q8fdAzwzdtF3w8/aXvAGlc6DfSFX+4uBwWnnAiUxUMy
qqqvo2iog4RiNwJMBceRVILOHx5iW66WAIdFzH8IbfiI8jzwHWBuYcpICa4Tv84UW7HfbXqmNkgF
WAiGzmtkRCoYgb8gHPTVM4HkjDagxKJzFpfkgDTFn7Cul4ScdhKfG3+V+o6gCSFdBOszxwRbGEb4
WbKncLzUEvNILwUkxYqJG3QqAqTBllICEo7MWWvKhB0vvxn4bEYALMWa/vjVotpc8HJviW/DPppa
UCaaC/ZSrY76+cK9qDvvvIGEd+9G8zr+s2KfEmE58zDF02tPI4Y3O8mI1WYs55dCxbz5PS0YtZKC
mOZac+qLpLUuMTg0KGlrCGD7ZAylaZSyXoYKCVauhW34d/g+4sXrGJL4Nu44YOoVDxlBWz8Nm683
grdybRUyfUjnm3tcdZHsMX63NZ44aR3nJvmHpf+tZ/FUPrnztNU8KBIr7QotPDkBvlrPsoffakEd
7u8wtnYmyZKenJ3cA+0oq7E6qfJMDa4nGmDJ7w6XERcb3R6D7+TKXl9eTx7loNAVzxrNoxBfwmy2
7Bs4HQKk3t3PlOgcPumfZR+bppy+3VOWeEsAblj0daX4Jo3yAn7uD95OC/HWY/M97f2FYHnfyugn
e5wb6hgvHvztZEMEFTXaVoVlnZAT44ZcMEqAiq480sZBkzNvQTpYxzmi5/RHTkHdZynoiALB306g
/ZUmvntgxunV9PoD/CgX7lMTWfgn7+nz+kJI5gS3dBhCTEAcQ30qNqbtrilym9Hbh7nQhw0mkWQB
oTr723ZZ/Wkt493fppJxu/DaV+kq+Urzvtx4g5ON5bC24+pe8rzTYclwjkdCuDLLOhEGrNOk3Y/R
Qay5IAbsBejZCRlRpdQWz5gr+Cyse/4NBgZGY8VUm0vfFtuCP/MyEtuxuo27S/ujJm9kH8ATEXQ2
LUbxuwD4ZS0CAtW1+AfMKaf+huO+7HUl5St1WmjFW6TevvljHp4oVg+TkOKDPpuRhgPPl5nsxpPo
5Kss3LegiYeq7rK432dTJh1cwhujxHOstxEeV30igHfrrc+jw/MfDeRcoQ0LCMByzEkpAA0pxrbd
212tTPP4oAfLJqwb29LneCQiTyI8+uKvaukJViaOSxu1nrx+H2JORTY6/KpunZWhrK7AKoVSxa01
gxhieWr+Ro2VjOfPdDXTPpdgRvkgq+1udkzBjlsA5z+zIU9/PVPAbXGvKUO1hd3+Og7xCFDlaEwY
lqsYDrbzBc243fm4yeuh+GAgkmXzL1BFeTWJQSuff8zjRbH6kzs/ltlTE3F/zbWVbo7Or+yyRnli
OwHfxDCeTq9j9NbgwN+8eehRJO4CYj833eHX1SQYDf0qnMlrRwU+zdHbOxJ8Ebpaa9Zy4+vOsY+8
IkH1thKLeC7k1o/SQrC0cmRJL3oLmmOjevZReUBvJc01DPD+zBjBlKcWdP2wLOo6nqBg3d2WkPEd
Whri9ZAhPCu2LsQlpVOLHKEiRZ74YoYzWpiNH5ERpXNfAHSrZjLs0UTEjo9WokCQRjNcpgeeyZL9
HlOZHHBDCHaVsDJ7AGH5QPie8TVEExZcCPMiTHLYfjJX1w4V5L5LlMZdV6mFOPsgSmH1Ddg9sWlA
aG23pSHOlTyGu2jK/n/xFWY0lzIoSzruBwwVaVZN9oVfl1ssNnAkBiOS9UULaJxMAZfINXJrOEiv
UmfvhQdjT5S2MOdjqxUHu6bwckYrDqx65C7WBURToZWd9gQWr/+3fpNOKtnfNEvpwxnoFC8/kaxh
juH4hAXLJAlhVUbafUWpgBI5+oqJaxwnO0VGhuiNu3FOGPGWjLl00IjGf5JyWQfD/PfZr06I8c8d
piGT1ylZ57gw5qIYZBs/792sB3PTkcsRjsmdXcM4LWzCv12u6+XsCJmfVdHIA0c6lpLy0CKRZJsK
9W9Q319B1vdrsBdqZHta5XJoQazgeOP/XHin0Izmki+Z/xynHsi+ReDkXK5VDup9Yo0YdleKVX4O
DCLKuFfZXHZpRy/goO/pCcXUChU3eAeWrlPx6ulELUiK8SNzxz2zSkaA1/pOke7g/IJbhUKmEpMU
0D+nxXoifdarVZzbTLQTyGJmlZfqNka2sDMYMAlDlOIr3uRVfTYX9Ve9AE4nJlCyr4AGGjHjne8Z
j2mrsvex5mPp2KbpUbcOalICvJXBVUau3Zkpc5xvqJewm2c7Zhu8nrQS9JAX+wQRvM6bBmW89Av7
8syvodsNNW6HAner6EPWmg0e948xKttmfYSpg7PVnd7CgjCa4wzIIze5vBbF5raMsql+LgMdmt9D
UKXVNTs0W1GAhFiHjJixYW13Zo1+1EPGWzjY1f6bKpIsU1vqOPDWU4gU5Ee/0c0gniY/drZz5k4b
qr7X/Y+mmiHPoNwukC2JIhl6Ko2amAapXjFxNw7iYRfOuHiGK/av6fxwGvzmHW0UPN7TJxR2Gh+0
UtEi8FuWUPU5WokBe6RB+/iIE54M+21bKQP7S2YmHQk/cvfVtqFihzMw8RZVq0D4yOSbIAu9g27E
qV4RkH+HDeUhjNqqelZiUwRRN5TXWPOBfXv49iOYFNhBsOYy6lsQIFX5hWzw+a8rOsvXIC457a+C
3QKi6g9hMtw88BzJI/2GBQwA48nUsmVOT2kLEBAdgUBDup8lRpYqaiAuxPypZiqFQxP2qD3RDp95
1Udhj/c0qcyJXP5Kznr6dI6Mp1yYkx5r22drpGbZcaCxvaja/VZ4hZ1UyihY1IZhQRbTi30jyT8Q
ar/OgpFyYFtDpQacG1UhoHjv3nXKNHX+4KRVIi1XsTSw5vpSW0xAV+T4wQLsLEC3UjE8sjDN3yNP
BK4i4xL3v2mEvBceccaXPxAnDCFhfA7q7vRTa1utQQ2IITeuN7twMlvNY/RqdXqJzOqheGy6SaiO
qumOhyIK5hNytFTg7idngthkFeFzufgjHmsgPhN4MMM6Uu8cTyr3G7ILHC7C7P/rfFcTN7bfJCBZ
eWzyVo4zp3w5+X1IQuqgROfzk3TV4FzbreUoq+G23D55VoJUux9uQSJiA9sRd3Rmw9QwAgC2Ehwn
QfKO8fM/bRH6CObwI/yYivKuPZW35IPoev4Wq/gBjYmpLfua+v9BnkiMEYB/u+/ZX6YVWObnw0kg
i8Ay5VlHRhHsSizvyCj75wSR8KKTFo0YSnRGtrX9IGRDTr3aI+OAjjj4ohDIKcfxmgOvSycygZT3
dhMAlgJujJ10LSVKjlk/SjWzN7ibiOqf3DVYnkXUprMTQJ7yrqreIHATgeckwk9lJsmzB8Z7QFCG
NHFsS/cuVIvsNZsEG1lIOmZ24gnpo4eEe29RFE6w5dlJdMS+pf4xoo0LM+nRVgj8Zma5cAv8gnu8
X3veaXDPqyo7rMsY8oehHJAkey7/oHebkv7tjAz/QdV8dXfN1m4G8GyRNRVkxwTWuPYRcAg4/8X3
YRCJmZmERa6/F5XSnDsoDsZAs2RdyVvMPDtiTvqRqlET+9slr4aMFYDw6f2BAIAjgMKOwrdIPL7Q
rYJ4eYk3rbLQd8gcidvCf+UQ24xO7LoN6SM8odkjRGbo+by5FGDKVmm1zyvZO1vDzBjLaju9c4xg
PSoz8q3rHnY90FGUOIVvcJyZ5ZSMLPO9xO+pW5RFZyN1QzAjqy/uX4aMYeit/d+Fxt9kSJ0venCd
bVcWLFb4NLNp9KHGFJeDPakcLKzEQINYVqyWlIqPM2xonHKtHakc8+qpjITX6mo/I/zZ3b2MqoLa
uMj7uqwtVjC6MsyJfnF6mNWWrm5jL+77NKN2a9CzmQGT9rkPj+tnBkZEp0mj9rsn4fe/JR34d5Iy
91/hrKooG/a5Tg3brc8On0t0am5m3zXc/dyZurZSIgHBL9L/YNIKGiphe8O0D3lVFKl0Xa8lAUJ9
JNfIYO0BcHeGyG6JMj1CLmMF7Mihp70eE68B9GgvIR7umbeVeJ+RHghNjPHfKVHmvUCQXwFGUmYN
Ur+fwkvlrtTAB5E7hn9aWItl/DSKxB85rVIiG5QpCg7NTor9QdLK6jecHoz90Psb8inT0ek7uEm9
6baRe+ZeNmV9eqYmCbz52uLOHB78zsoobH+cEV4qroSB9kXkN4O0bDEEpaXTmOFzX+/B2W0BCz37
n6lth5tX8ZId9ISjkdib0mk3r18RllOuynp+DBv79PTsoM1NGLEBPgC87ZKTb+eeSM4d1dWiysc/
Wa8805oMcP3CEQWAKJ6Lw3nLWylUufERvCSckDtZxBCRjjF5Pujmbr6fVk+I8JlPfrDzxxyHkWgD
0Fx+A9bAZiVXXTl0KDVyVczqkXv1Hx4Q882S/QSgl8phLUXrlgfHBrSqW5XCd54a++8Ss7W2izPL
a4QHqeOlJ27XA4D0VylY4E0SBLu0hYdRZ993mQ8SydTOGvrCsLBVewJFvVx0y+gcsa8yg3MXTea+
DtFwQPiHgVjFBZJCB2Owg9thxxlEV2IYedCJQ+SI/vHsAPxl/k9OrT1SYJ65Df/3fVhYfSWPPxDr
BY+Z+WP7aj5Ze6K95+ZUl+l32v0mgU3WSOPvHJfGwUT0D66C0xolVHRNb+KLiy/5zDnuVR+8qWkq
yjTRtrXLrmbVH18ixWriHReGFSwkdsf9lDcqrDEKaMc1URYfgeqmVGZZOAxKl9V/DyunR2oZiMTu
IscQGWhIvdnOsbk//7dFQqPrFblHtlCgmjAhfQFCJ8rFP/HhkXThkd/OvKQ5jjzb4B4Z9ANB8dWk
Jiwxgio6HNrwyR0lf+ATibINliCxveYfEgU/feHVddc0EqMuUnO4U6Jk3xEuqeJaBymd9TrCRdJm
jIwhAf2JvqOlumK8UtlZnxpLbABmrOqH4aD2td0oy6Ckkm8ntuA4RVUWUW0A3kpXE+PoFwaXLXBT
1quZO2o4fqmZxiDXR9kEE8tqz24b4tiFadfzZ63DhEr+23P7nixJhd6U6NVvDDoTyHhJhzR7MMKo
8cX8dYqhRkmaSfKJh+KPSXE0a5AgtzRqcILJIxJe2tTv+8EVV+OTSls6RDJ6Udnf1lexzpu8H32R
IpvdbichwfUJFlJ/7ylZBuFBYBT0EpPZ4DaW7ceVWgR84gzSyvMhrQbFU6+Dv3dT8giy8r7nMD7G
Gv+ATP/It8cYixIAKw+kjZIzfeIhwybDbhOhaLVkWX4s/A87GDKQ0I7cHEB6ilrztSv1jQVDiFLP
qSsPdo/eqfYTu0NigBr4rBsOWKAaFDmOf97Vx98Uid2AYho3HEieBjpP0sRnWdmtdRSBNxzc8V6f
p7T9MxKH9jRnbbhqR2HpPDBs/22bqC6+tU5paaG6MGpVMMUZjA03luDCu7lsBxOwlhUNzLYtxhY3
a0P1qyZNmIV1dXCrzRuNrA79jQPlhZ6gBEjVDx7bEu67JXVDUdU1Th8E4ewDHL2wNHbVHSgDTqM7
3QYiCvD7RVJ+jWagdfh3gtlHtSaElegQ2Ea8H+QY6GfCfqfjKcRcIsVTKz0CrfRs+EXVr3BCRl35
3OKOx16GUxpy+9oqnoj/RaYu8k6VyWoScc8Ih1AlvFFDwBdCtLMjnQJb0AzVVcdJrGzYV0eqIU7x
e9gvl3xLviAdcdEYJhlwuzWSAHwLI9lrGhgF6pWcCzRZ5BnpGkzECrvzlyToZWaqAnJ/4cXCpQzt
H/V5q61Caqt7WlVIgJ65npVYY0DUq16WhpX5vzt7LcXzszM2nWnWCksV0waei6HZlf2lToUsVVla
dQKZBwmZo2RUEMUbAAZA60FeStWZ4PD1RyUrQfmav8TkylsJjRbZq4jtCS/xrGzHH7C6Ex5nysRu
csU3VVifxTRMb8aUwLggZkObGVrjyabd2EUvprvRcSbASNUwtMr40pnnmuHHVkR5uT6+oov65+8S
pYf24/IaZd/71THgn7Vk19KGGxImAyVe1UjAhGEEcuwjzfZzL8Ri4/M9AtDBlO3+0q63H7UQowxf
16RJ74MDcoWkjU4d4R908+b6GiB+WHqxeWT1ewRZ4RybzNGMSIPX9B51Ek/D2NVJeehOA6dOZPJ4
LXQbnvLMZqmqBPNQyG+jWDwMHogUcsnXJosC9sf8O673OnVwG37jJsSHKidnamONDsU5wydIvTIY
0HIG0YQLC2sWP++SneLD3Twr8VvQ1e3LTPfldTOvp9RhjGz1Mw1aUaIOJVv/ANq3Dw/26Dhzhvs0
jpV/5bDR2ZuDBv8V50kXpBs4BD/CFOxnj8MDEJrUZ6ke5Cm4puy5yxbfDcqfpVJZeBTQOWJsTjXu
htjSLb9V9FXp4X0NFgMNFKgFaD40dq+k8QCucqdWZmQggUdnlJMDfkklekPy9z/kp5WRbTBeEbkN
38U3tOnWs4zallUU0EcrlDvO/zjZ+dRL23XoaZunB1A/sDxXvw2F+M0gV799ahjivadWSuJp/1yS
lmJj138hiZyEl/ELdFa808Kz8PY4hn1/ZSYkl7UZou8TzZ2GEuw9tVplY97Coc2qK45w9wzISIHn
xmFflD0JkIXx120+vl9I5gDW2EQz/3KhUy9FCze7vxigCErSRFq6HnmJiWYc1QL40/x0p0wNXUvI
laZZQAfjZi0embGZWuc0un4Uxu5Q7U3h2V+1L/Q9tksW6ZI7uTHYRw4spcH0HfgoupCXLoYmDuiJ
CKMUQtJ+2nbG10DGYcYXX/wbEo+pL95EdV6x4beJY2mbe6oiSWNFwQQN37V73xs3+Mo7EFVlG1mP
9ocZWmK29wMnKy87DWUc/SGk+Do2BkwTXHz5WP3NTTCKMfHcYRvY6A9ngqD3UwXF3PtoKq1k+suS
ZK9SGJTd7L0vXM8CWaPWhHkOBT2wOTucPrNpWlcijqS015QABccQQQuiVJMRJEj7GBBlYgylmlJm
AU5UX7a32NNv2aXUjDLAYNceX4XwiN+RwtpA6C8ghy/25+9zuJRIlUmwdXJUUuI+G7o5RegjfrqE
i+JfpQzh1l/Xx6NXyQuSQh1PGClk3fuSR89nacrVdn985qsQBb1rHsHGPJrMFCSQT++wnO+33tyl
UuE23qz74zwL/LmsghnyAx5798tNi5IODBNW441IRnKdjow39pdWqwGCVkcITDcFOrUgRLtVBwwp
q4Rl7ewBw9CKBEyt3r33XynTGmUbIyByvlwkpLaGm5s4UcUwfwkIR20sCbJJhbwIE9qJGbNh7+Q4
Sr99bdsDTqRGNZSX2OcH4hLNt1WhCkG5zBRLkhD6ahri2WGyUDZtfi8OXdYWR9pRBtY+AHKF8Hob
wIB6lUzsFf17rH+7XIMju1/FPLSFIr4a77t/V5sbcP+qKEfiR51ycQTYj1r1xSLRQ19ZR1+qxkfk
fyoMzrrVQGB+Ghy9t3yJsLmh2ZyCEErba3sQOZfh3U8A87JgxPN8vCKDrV/yGHuiNsZdaAoDb+9G
E3eBgjpjhzCcmYL/5zM4KGfogLzZD5zAetkoPTiPAWGIupNlqKEZJHWXtP3gQ5T1qkEZ/9PDnEOt
lidjOExeB0DUA2Hask363xJLBeCBtewbu790YrilvNW+Cnzoc/HalBkzvtJKM97BfcoJxr4YM7ET
oPVkCRwPlN84ts+RJTYnKFFedr+LkayUMja9gB+XNEZ76OXAs0JCVNLHnsBfcLjp0+UGIdAzpH6h
IYgSVOF980vWBGp6Yn5VjjS58xC0Y6dtYj32BjR1QKmsspsg3MzATPt/dabf/eS28ahFFBpJfCYk
BLb87Dh3jOxOU9IGIw1gvM7S6Zqml6k7H3qyYyp3VZBIvrjpg5pdW0UUcMyVf6cNQt+PShcqC4Nf
XFQlFleLEidVOln5fP5NkyJzaZ/+abVsnH2+agg02TTn1IbJ8A0w9bn5s0s7RKrhMeswxDx/JDwo
iXDpFEqIegHwD5JPUXZvOLNgepjPLseCY3Ce/mt1FYZn+lst9wPm2sT13roYVohiGg1qZF5mzVqw
cswv7WYpjZp6DsRMWhxKHHqfczE2lWwbQrpyYj9Lwsbb2wVrBaCuqDBi4gQ78vDTSR0Aq7UnWbO2
4Uft5HEpAVMbwXy1ouFF2xV21czJDWxBjkjuIiy/fb0CoR/R9ktze7WxrvoewTgTp/TOsqQtRzQt
rMIUrLcS9clTl507PN7Z94RPAZfZP/q+c9+IMXhHUOTyHvE2o+8FD9Hmw2v9sOuUi6TcOcz+uLhN
Mu33JLPAlOSJHPJSt7eqXxjr7krsXvL9BvWI1gbYyEUiUFNIGbOf8xbGNgLIcERhX0OZjRPdv5jZ
HCaGqnddi5juL32ARYSlTknKWK2rlL2RKkipJVqeA/QUrRSI8doTfxKEOSDFCduTMERfqtAaoCHu
sv728qIXMW0bVLTqsNS1bppAGttI2l6wEz8RxQyogdsJGgX/Yp0N1KvLVFLm+LcHok2HTCJjfQOc
Hu+S0kGapfiikf1Zy9ZKvYlyJXe0l1zauxQSqJ2hjbGa+fExubLFUgz4UyjH3Dxrp9m+QfXtTzIl
oyZk4BETF2VxpaBzj/Ue7bvZplu0FB6FykcLYDhqs4P6HPVSfz4Yio+mDwXd7oO/r8FLD9eliFJq
HeQjBQQxP8pjZ+HkQb9hCrwCdaeHySnN1lLc5AKhhbjA46FM4ALd/ffZROu0qPrpFKB7KyBcpSrA
B3kLArPMtUS2GnL6Qf8kvrA0sUHf3CpC9dec0t/On43WoaMmkSChvyg4JSoAIvpL/6Y6cuCJV84R
axl8TZf9NOJ1AXcaA72iloBrSIdWQZzpQZi1Vxxu+K02bsckp5SBym2j2vunuMKc4GDNVsLSRO8A
I5JNDLXUNGQG0U2d0p0o73dunO5cj4yq/B9IvpgT4NPVaeRMMlForBQucAU9FrETGaERWCe4dR76
LtNEweXfyeZrdz6qAre3uZFxRLWltod1jVHO0hMx2H7fLYivK+X0rkqwz7aZ5CEhuEzXRDFJunIa
GAH859BS3vzijgWxv1D2nvbiNVyKsgf/+chn17CDUKvbNneHqk1zOLhLbKVaW9Lb0QGY/DsZ6Mct
ysuxUb0Vr+oFA85aHHytJVYeIOVanlkHjXICodUnquB92jVfgaT8lIiuJ1zxfjvTMlUZMsQV+PpH
FqLr0ao8ODWug3kWqgPqmk3C5y0g8OxeLmptx8yFCbZNTf6OEWr73TyUNtnG3FQwwVZ+aeM9HuKE
RwI6YYyiZNpWpB9h4FFhe96z8ESOOQqYz9LO6CcchnYzKkq1Etjs2Q1vpTClAqRLB1VLTJ1lT5GV
jK6l0nWdzbAwaygBfHBeCnnW9ehh9U3eoekEkuhKQaiT616KVEYSpCFoAC+tRKEq0Kc+SS7YqeRv
Ts7enNiNP8J7zrUgDjF+MogIbJ75Mze0kATL+l+MI1SMZIlb87wHoB7GW9P4kN9Fd6ZnkxQre0YK
j3eGqEyTdf+PRIHr/VzTt7boWbglaElCah/QYdTWAR0rRb+1z78nBpfxofv++tT9qLuVXF+nFaJJ
HuokvzsJuZst/G5dug8ACp8gIU+Lb9tW0aWvwwvMZ3pjDq/wOnIotRpVhV/qKj2FbyFvRzL3d6HP
TOenImyfvZJIW8aLG88Llfer07m+X6jyuOmdb084wtDT1ShI1uMsdMMiqr+9Rdqg1zWAUDiFXZZe
+J8NknB1ZSncAr17w10YTbOXezCcUV8Ge0YYgShMXAfYE62v7yR5sx67lVqotPWHiHNNkGD3vxnA
jTCL83qBwJrjp+Vxv9kAEFBsp+zSKId2vtmt80aOXthtlaoY5TzAF9zm/u62Hfl2Hv9mlJBD9/XC
II7HRFJCSRi5X4s9uoSnXB8C488ouh992252WfDkmhup5wQnCQc5S2WxuySnBwKunyMVyVxy6y+v
vjplreJkTFQOEu5p7v12EdGPxTn3p6aFdpxkeaXqPM/3iPSknNcqK8T4jxKKvYuGlyQ/m186iCGb
oOZqadNxVY8pRUv5rIU1pHPk7acMFEJZHef30YxeftzEdikVP8xX6cq9B+zxmTpMOsY9zV3cZoaZ
Seb5+fr/r1sRjB8baJVig/WcYCPDc0xnggmaJ0uEGZKkwwXjWt7ggwI0XO+nSq4HGmDbQOnl0748
HptEHEIVwAhnLRu0WusaHxVHcmr+bnLLl0PwOodeRoqbw93P/zwHVQd04pdxAdz4GXhjtJ2R4aNN
wQrwMiW+0CUkWSnhXLioRhuonJC3lW9eQ5A9a2uSiqaUgm/brDt/oaQaHazhwY4YoFsq0p0OCyly
Gmv9BKJPC0UPsucyvCRinuxC48l5btzX9DeR18IEBvfa/IUnEO0Hj0cACpxTyHBJJeDC34HbqM6S
0Nh2GRKqSjA7luyNO1vip8K/dO/OnsflJh8qar0E676bNvkSyu1/lRRAuq8lQTEbSNxT3R8R4M+x
nmQ+CYtvZmxqLZQJxClp9xs5My/Ki9H9de4WTyMF/qalWBGZG1qW61ANUKkGc9aH0cId/Jrslvdn
d9CXrDLbM/mI2CEQCN0bHeYuHZHTaGbhV03TPv5Elk1DugCkdp1ptPIBA19GyJBUonljY08wBjJC
L+nxK/7MzTGV8Ou0UcOByhH9/i97XY3AVA1eXQKs9Ob3nbP3ZWQV8hD35z5XCvCvyozkb7LIqavC
LC84MzZR44NT9bXBBCv9X6RzJxXF/uqxGJ0Ip4g9LTA3Cr1+WJiaVybBFGIW4vFwUgvEvVuQd8Bk
h5sa6DlTidE7WYzZqyuMlMR7Wtc+jpZUKh/18YzX9UN4aEdoQLbuvT0lzDPcZUsTvk0TniI76Q3B
wH+hL/VcfR3iDWvQC9INMx9fr7UO23D5nt0RnyO9vBzCcKrTOcUObw/kLIMVdYMKCjTUvS7/6b//
4z2Hv8MUErbwb6mw7TMqgwOvwpANLcLCJvOanb6Bdh6rQSlTkpD9z9/xVlYSEP0TFkLsb71AtwC7
jpaeAM/ijy2V3IaPIWl3W8qsXHREoIHcMWnZG12uUob63kYOzC5kAvmpAX3oIZOuw5PQG/cjUaxs
x+SsXoUy0QAt6CwOG44+1z/fuFopRsf3Q7ftyIXXqnehAR+et54upU67ExyKg6e6Zbh96DOShM+c
ATeS6Qo9TU1ZEvBcbxxd5doT/ZiOwPzjT/T+riCOh28viMrJPT6VhXC1wfOfv3vA5toEze+d/a30
j5CPcPyQ9vCigRBX9AxA0h/wxDqGhtvVCglqypiE6m2vhU/sHWD2Y4exCleLtHazgyCTAesc62Z/
J3l80gNGgf/JxAxM+V3XRc1KuJz9ZY3mVbshX2nK3RO+8IN7Kb0GSgvEasKqh6ps1TZOPcncktI3
yewjbxxTSHX6dOQ0H1NIUXUaYu2ybNe+Qs46zql6cbGt8pajjQF3X63AzyUI2MkffXyPPcqZP1ve
MAYHh+RFBSdUSIU4ofPRSMlG6wYhkOZB7d1ZJ57eFp4fVbiSIqU6q/31FWD+VlyGq+D7OsixdJdd
abHp/CSnIkJP2nxAnZK3gHVZJKBCbbSJW/S4N8jh8v39vNjywE0w/V6FzXsPTNPwfTEzVvvWJBa7
HjqXPrNPRfeFa5WlR6wsixxjFIjcnj5Cksw6NMXsX4JNtRWTEwtB8rgnLnYpCKsMNGBXntABbu75
qkq2u8Qo7OLWBI2o6ojJOpKI+RnllduD2cAqM+rQTF61mpPoGjt67K18H740cTXysww/QNKkxqPS
/Yjkcsh2aDJZmPVZ+hX6O5+lV77xT+vWSK1i3sHmrof1Kkl8J19qbsACaRvqH/DiB3oYXhFEp7/k
OdTqrjaaFYSmTEDB3aAjVHVDvaKfojhuJLn6dXZAVC6a0HYLjD2FAHYMz9/PsMFDOiszqar9AE7U
7rmzNsvCpCIC8mXy497cJFRUy3Gdw4DV2zymv+HIJ14GCi1tKY7Nxq9XR13rESqaKwBnwmyW0jUP
KFpoWmFJ5MCTEzWBCPydM98W9sE+ztpQzSUDn8eiuo13u0aqEAY1+VjEpCR70B3r7nHsqYbW0Fls
UMUMmkR3GPl3NFayebzjZBr6xrN9fwXBbiHEF/kyrOUTU4A0BXowBZ9k6f45qYzNSn9UrXoqrBDe
BZ4N2Nuiv6tAd8xkOXF2tUwbVWfcAJxCc4RAsWIYmmLxX3MX28g75uVQOquRwkn0XhxD/3TerFyn
+AR8fnCLrp7nQAQia10vV5RFKu+MhqPL6L9v/zDI1AigZD859kYsBqWWWFAyAJ0NYyS8hKhbVfpO
S+vBnDPJDl9kVlTuic6qYWelV7jduFmtDoY2vc9XT8TKJQG+bHJOFPI56qG3MRSfZuQmZYnRj6Ch
SOhnGemivcbkN/qPMjbsDw4H07bYoVICWKIq+SM7llIv2CC4s+5B21I8bLczVOLAaGxxY7ye3IdX
hIOaiqhr1Lz/XaP6y8draNBVLTACshOAHvXxNrGYCmIQ5eNdSxFSfXgQaxL3j/c98X/n9COuurBP
09zej3BJQUtfb/8zCtUbGYKD1YTqGsH3AY2vPujoqXCPERDnGFzMU43rAnQUWYCkrmli1j1ogyXa
nytUK3CgpIweQBthHki5SNPVAj98vXSPSfz3EKw6lZlIXba6KlwjG/iFFWNYHLq7zapHihYKX8i4
UN0nVm7B0yEAmvMRIE9lrU07iVHB5FalLYFRAEzRwJD+TVKQ2SvDQJiIQupOiMTIzdBBVfhBUZXW
AzmrkSUDgbbFtEClch7ejiKFpRxnuD5IKEbeyOSELDy35ay9nXJiU/xH/hvQBYQ8MDXtKdRhsnFb
McEY+sILI/d+zVB7qeeh37suPalAdt8UyvZsDDxQpzexOCMkFVKMO7WJabzcolaIy9exc/GIxLiY
DjeBjLS13eWNE2ObZMgI6JfIFfaz/3z+ZWmo4RV+YltO2uZ1zpffUfq2jpgAt7eaqv1ppmS6gHZ+
HHYiMMXh4TAAvOD5wMIK0xO36QFHVrx0BMsIG9XPBYbTOW1rrol05yOnjmJ/zdyPVnmvSCizbKC4
/7RtCnw0Y2wAqwxYCrNRGASbon9WVKRQ/5/zLibDBBQjht3s7vY3yaCw9nJiMSuNR8w4PUEHw5f1
27A3QpknaBYHabpOpQFMlWiSQcpv+LlVnUn7FQoQhRADOCPKdG95Y6F/A5Z1V7N+5uBwesKoxPf0
V1sSx9tEAAeKVgOA+ZPd8aALhcnU6ShBn4L4CCppotpkYPbMhqSkEl2liVqIniSKHKKu/ikODUhb
+UcnLsKOGW6SUHZwt4G5NAiv3A61CIsGQXbvZW8FCuQt84wcVNdWR8d1j6NFjUg1z09yXjGjeH4D
6t/R63qJI9rYgVuSabH7yusmaDmgQ6e9zo4I2nXWoDy3Mrlhk7flfyOBf2wgB5k6MuZ9gH/i5HFP
HSjJe5gbKhrYLMKQXSUdkTI2JZbWRQawSWIF8VyPlEEtga8mhKs1NdYjSlRgA2HXxtlS30XwcpGb
4QawtwxndXmPmVynXif+jHGUJoDqBaexFyAMOGVVwnTY7OiqCpus46bGLjkPMMgzszDZHU0gpAsd
4BarvUDDja9VnXfXe4MMyHcOLh5WNzNc2PaObbSGnGcaiRcT/goGvcePSZKJElyDwFcwPL/Wpogv
s4YEXWdGRrHqAYTDk7L6ps4k3LoajT7tdzGmk4+7nzaIci8aR0KZN0ibbCJU5Bb/MAajVtV/Wb6g
lvGMdJZS6aIeTwBBQoKOsHfhamgp0qeRZc7M2SRHjvY0NgQ312zNjWHmIZBSiXL/L7KlNC2Snidg
36Z4RB+LS1zAZNHlV7zmjdIQGlKjiE5njqlAhNvLM8fbsNkerdr7mZHi77XcdHqtxVoIB/rGGMCG
k8UGLLbttpCcpo0SgOTyujeaUKCozAV8dhoROjsFCOrfBIJw67H0ZXtlBHVP2NuZvGjgu9TiyMcQ
Qwb9PI/H8RIIgEzXopfPZCeW+1mQ8slOtpaeJAXI3+A+8mDzpNMxMkIEKdM2NwskxQ3Fc5sWlLhS
MTM1Ma1qgQuJzZAXy8di2A426+tsB4s9UX1uHfwCUDZYxC1qvkjH9zi7yopSBBvyEzIb2kDzBqdm
Dcnm1nsU/b5MC2dHGryL9+5kLUkwMuZ3vY6THIs3RjCOBZEjzvotuPt0JF2v6QILAZl/rrrkpXTS
yom2U3U5Q09afDpdYLFulG/vzjVgvmOkAD+ovNWOCGLg9kBbfUtwgxOJBkm67SBMZNUZ6Afb4ZzT
YVEQfj4rYHqLMaJ1t9jhdKlnKVlob20Ega5L5RGMApDg3O7M8biF20xNTPLqyb+PkuAnv0Fr5KHM
J1vzG1alR+4cSIYPv03aB+pC9fnogQOyq/xLv5pPPU9fJZc60z6XCYuW0NxS7eLGv2s92eQ8Lcrz
+h0dkMvEc58wMlJT3CSSC4KxMt8QLjYARvBeO27Miaz4LqsFGYNbE5JlbIkHWliDYT+m+4cRJACc
KNJwsV9ewkdciPrXoXJdCCzBfE15+2aM3umAVBYa1COzfxC3tm1WWAJN0PadL0fkyyFrI45oSalR
Ft8+QKsXqJHC/yuzX86WHzZSOEzoffV6Ga2Ef4aF+KuhebXGVfIR4qvacst6L8xB5JH/44QwrFS1
FmMNFSU0fJWC9cARrH0zuB/oULt09DhV0APE9VqX+pn/w3eyI7T8eDpERG6J6QdMdMKzkmQxNAgh
SD7qUklAKxss3T7bWhuAjjKO5z8g0872GFK5fuC3S3QMfsB3kGpX7AyAT3Y6+A5zaEb0bunZLieQ
+FY3ifqTt8IpJXYu79g6lHgDjQngeeGhQ/oW7JTeN7fiuVGLAUO5HNwP+eWmrp213b0E5RlgVRnJ
3Mqx91nM9ufJMAizyrsDtWNLoM2lda9kYQNnM29l39ibIzf7bnNurSrjPAqKaVeH0uUMGYX+NpuW
oUXdHexHvwqyrUAU7POy1GEWUUsb529Br+JF+IgAvhJ5dFcQ0uheerCeBnXyH/Yk4biLYemkpuGG
fVTsnuCX93ckHci/DeBR6euTMnFTu7Uc4ZglV3dU1eapuA7u+pgZaOyq+5yZlSxoCjbIdQiHMCnv
jkGjBOHAbdSMnSQ70ttbTiim7/HDQR5oCtz+7sRwPukO/Vpb8SRgsCzSAG4HyZXhnAtNrNATu/E5
efOvKVFzkLW1R1Gad/ifKwQhLVRsnDb1oC+VjhbucNidcXsFBKCwBL0SVbdYVhLccj+owfezSUBq
oHW7GIc2UJSIe9x1sco5NIXxRP61GaNfgi6099Ur2Ktioy2bjxR0KOyHZSf5vgvu50kbl42jvmAF
rzNRHyBiqNirCdGRFD0JSIAat28XLhwxiDWGFd55m+J5BSgGo7KgxUavREltQdg3fcuxHdySizWK
W7g6Kp+H906UkOBc61JVAQTZzjGDaHiWk+myyrlNChntOR/KHBiEl3BAH08na77J/J9B9joYIdkJ
lA5owTRsCGhX91XzAFNZRw2UVvO5d+IqbFlVzb5w1CCCFFUpMUgu4lf7Wx7rp4r6+pX1umW9vJ2P
41TmQ5wjih8qYJDzPoqxXMj/UVmouHkXYXxYe08TTXrsDJZTwBdFm9lVpu9pJ0b6CDAcvQ07n/Yf
6a7jrmy9+fXeFF90Cl5wUFRXTYL5wRa/RSIGIzjMob9EjtgOJDkgHNhY1pjtIM4W7noQxbg2QOnE
1ZYtFX0H7Sgj+rL1qc/sSPP4HSFWhK21k8dhIkTU0MQvI5FXVNQf8Yl9gWbYFyyL5eo/TuDrLGSr
ZCG4zPeBTgOjlFOb+goNQExNs4cI2E+yZAjtX0I1bAo4zhsAcTAIv6hKlwKijHO72aSEgYcakdKV
QMFHz1RwupKAgsI07iz0adO4wIu0uxBJ3/UgsfcGXeQ3OWIZ9ikT3JJkGiwLBZajPnz/rR4b9CMF
ymcUNKKC0G3HSvnUSRZmUfKodwNEIwlhpKSpfKt+TALxC0vuQJZzqEa2amcYgR8ZY/8VfjStbvXq
/BOZboc8CWSRvZ6sMQwP02FfcLlzqS6+pj64FdJbhLu54NyeQp7naq6g/vNagE2oXOfCnbF48tWN
SMKFSrQNx/ugk9jEo3wMV6hyC6Cc512kppHt8R6m0388EPf1I6ItcQRWQpkLV6tNnbldhM0c2bIc
khWnj+eArm8EneXsyHIZwU75VdeQ/SO6ypQnHRSCd834ta+sdVFsp84nHsZoB2+VTLd+sQ/ar8HV
uGTTlTFyec36zRK3It0DDkcULW/HZzPQcouS7vj4tSf3letB5KK1XLB62/tbEkSBv5XvgMdFw74W
60mFH9K3kGauFbqm50Y88sChXujwmZHbkLfrS7oIeFpKRBbfjCgrXPZjhxbcmBk9/z/1ZcuGpsnW
zLT5qeYQgSOQybE6ULWK5GhVRtsRgHxasfdqEqNGOWiI7VWhP+1XwSIWWR8fFYnLBMvBITsXWnhV
0QUctQ29oLaY6lhbl/6HoSKVOEcO9xneoPhvtdOQ+LmiCWYj9W9szFI9Kp7l8f7ac+lQoeiFLdzD
rBtKvhGLkc0omd3TKhF0R6g1wG4MwZ914Q4O6fkmcsQotTxahG2LWw5V/4+a71H56IRDwAGfYzKe
mr4eYPukLkw7sBouzNBeOfkfjaM4myW+wI9r1gEaC1rQjLQEIC9XGwjCgkH8oKTZp57jNsOZJerS
wx4GfwEFdYqKh2cZZcycbNeax+d4+2bxZnPbGg5mXp+rz3aPXEGMz70k/ZuCk3R/JVyYF30Md3au
kBcNjC9446+smpsZ3D15v/ich2fWfqmdhGYj0HRVNzsLpy75Z2uIMjBvaEqXoB7FVsot/4D10c7E
g8IJ3WmlqJYDt1Qz9i1S5NBXzjp0/xdGyzi/W+2wS/LxtctMsbP+Lf5BEGxRGhWlJAw3Atwwzwmo
BLPtYLNUz3rfkL28Yvz4X2ggRajmmEfjWKdHUcvF8Bxz71kwU6pRT47NBoczqBsdIlycjwZiS72m
PjnH9I++MkISRCetayLYRH3RS0ut/YLHJpVRmHEE7u4B8w5Hvj4KWwc7coY4gYzOZMOHsamX2vtc
/30vlIwAGvBmjOl2U2DmpkieYfDJ8AvU1GRkexSZI5ioIr+xzoeoNS1tQ3ybGAvqFaG/LlDQNZ6w
a31W/YyaiVvst/9kjzfdRqpZ5wXthPfrvByqvCt1tYuOLra9Aoiq3KDMQ2d16+37UFSwMq0xVgGP
VpYR9xSpb2p01IAn/zN/lx25si2bLUzJI/OMJTuTRww+R01b+JlqcjKmtivqnAky4ViQ10beYFQT
Nrsplf022pdqTvnDj4xoq2esgVZfb+wrQ5yutxHkfWPSN37krJF2Gz6EfRxY68SiiAqQkdgJ2FN6
0c6tyLC9wxhD7vmktt37pzyfkrx8pv4z6ofQNfaJuEH7xlTmmVWwW1hITwzTyt7n/bsnNoW/Et1q
cJrePCTfwig6sR+szn/73BOO/ULs/GrPMz6GVsti/u8KRZLBWhLOXjdL6uhsewypXvgOkRJGEiMb
yP9nBkALrk+cSC7Q1j+g+oRXncAH+CsemUOPUb/SRNVp7nkiKX7qn/GxFXjJvcyKJYbmrDy6cjiB
ka91sXhetas7QJFHb1wi0B0gO1ym3B8aOyUldRtqZ6bUaOT41L9sgHhtKl1ZpzyfVSKXWEcPSZNm
EeDASUMjYWv9xExhI7Cy38pQn5Pu2/FIL1/ARcHi0JfQANiYjqU4CV8rSpf9+xXneanxckceiV/L
QicNEHz0mp7Ydm1J90aXxzv+eqEax2heztIQA5LMXDvE7R9oGvO7l4eIZIWTyUJsn2JhQPZUqcCs
f94zLeY5o2urOjAg8v9UViW+dhKZzLRMZlP0ekwVHV/RjAPI+8Uz1eCUEvaElST6Ub73J75OUQb1
6TqRLtJMVz9Kr5Bs/y3OFPF243BuDDXznK9sQS2Aqs+iQtz5kk4Phh7ZDt/FTNNe3YtEmQW7SOQM
38k5CLrCrRmbh+qe54DQeBYSn8VouBRewBqzjJky69BZ65qsvlNyOzygE+8TraZLv813+QC0XI9G
6RZBJWxUkALYTnmVKGc7O5VRD3zWZvO+th01sLsz/yGphxCyrzK/7z/etDNbfpPUt8AP3OdXkQuX
0c0C7T/VhTve9CGs/ok8hUqAIU8nzTvUMQGYEtTKYCkcuantonD3dnM6MXsplkh1AAb23AMkbXW5
YbKXofZBciYxX8CTwOUYZfdFhvieupdn8iVWHEKfd3mT3IP1k7ezmmzG3IX47c9WCyceTIxAZodE
zq4IMtzFcbNAViLZkq/CUFe+rQp+gnTt0Qx02VSQflsbzwJ2KltTwERcbFdKmer4E8/ABLgPHF5W
Lf0Caiih3BntWpyQ68VUqblXips6X4E8LZT57V6cRJFLPPX/8hFH547O7Z7aBmu4hDWHu9rIz+qi
xCjjrDlLFFWj0RR2GFXSHiTFQRrK579mGP5w+GAKZORCeyhAE19Utvn6YK94uKidatDBCpMx8pUW
FwhAQjN/8GQjUUgE+yETuhEwBxltxMj5cSkqva8qi/zR0TtReElrfvm5UlSl5rfgLZQaqEmrH7Rj
DWGgz35FIdi9aEWdXj2iO2z4w7j5T1f/fp2IjBD7bRHXahnCryqWPtIvyuSqkzKs7D6vWyfXIzYk
+yNbOC28YXuiO13vk1BmM44mwXumJ9u++LEFmiSYUhtI068Uo36C/3nZXE1YIlJlgyczCCfXRNP5
dTIkPGSEX0dxEWGs/gy7ZQVb5uf/U/q9rueJBVZPQyGoHkKN2+p10bC+nDRG92kr10dLpblOAj+n
d3u6dlz2zQuYllDL+VXct0R+qgn2iw85Nzr7fVR0EQWgetuqr8lZsEvyOrBqhl8nYd0gv6XVYhNC
w8VPRrO7/rNr1oub9cAKXYRd7sYJDu3oc0XbTLc5ngwzj1wVMTKdN5qINVhxolVtNowUgjP9ndKR
RoMrnZ1NvhBUzse7lQs+0K3LXvYgF+HeBFlF5hXONE1NuG+kc++dIqOkTPBKw7LA+CKk7KxoZWea
/IljQqm7U+BKYc2ew5zTSqIN+4AdN9z9G7n1S8X2GI2OppWlS6Y0rsc+HIVpiXuTfIzHImOs6ZE2
bsshFxM/o/VhIl2idpugeo7lolBkIgOyoK4nBSrOMjOrOZfJJz6otrRCMDFDdPK/+RiT4eAKAGqG
d/lUkn6qkhR41BT2s7HGW3DOPLDWCIE507fa9qJD09uIqmxsYv8BsTQznCMzRD7WIFldvHI44yN1
mE6au4LzfNT9ni33gzD81zVATa1Mk5ITDss4cX1IT5th+d+SabaCvOWDJSKTxmWhLARhEcyGNxzW
6QJIrgzFaTJLPWmdNi/cVb2Pau/ryKhLlvkGfvr3VUbdiYlUlz/i6gY5EGorMkfkYBI32lz6SUQJ
xHCg5I3p6dy3cvSLE85Cpa/RlPrrNJoD3rrdL6N+SKZexSHIe41CxIZaslEKXKwmgEevAPd6Tei9
9nIX+dMM73LYTxGvvAcsNrkbJIWkdIVdYYDC3Np8Ubyh/SCgOr/+P1QMYOSEfG9A82H5caxvCXGL
D7O/DtVEpBp+mUAAdDUxyydgbij3oOuyf+RJJNgCWjXh+QaMasWjvXZjFj5FRQFfRw9UYv+c+LvY
gBcoC27ixBTO3iYHFGOtxnQfv5bUpW94V+dIjtE0quTzNqEeSN2Ikm64u7ls2/TAlFuC98I0mMnZ
ZyOMI0T+lawyZwC2EzKlUfzJfC97xkHthVJuvQuGzxjr0DgY1sgADUsgU8EUpptN7Zx7rpZ5/9Wn
DRekiahtoUuEHhRLKqUKyNLfvq+inmFf6JqnWCkaoF52eCa9bYhcfvsy5suz+UruCVZKydQC7/MX
3OAr7aWsPEV7TUR1wy3kYwjSDOQdP95E32XhWWCZO5hh1tUp8HOtgffvzFYe7cVprxexZaD6wxS/
L2/O8eGIWcSkhBlVoyERZVvlDi9BNby2eUBblWgjjjJ2WSHa1P8UBhYliO4e/R08itvwrDnTaWRZ
9QY4a/ggQroT+Ijtodapxczl4OPZ05ma0T1rH1SU2t4SPQ5JS7URvczXOszvWpEr60JyJMOA37us
Zg6DAAAZpwLtkOxzd2WmF5+0Mw9SImr/731taYQ8PbkJNAoniyHDubJyhUBlbeeAfq9SnW818thE
UlpMtA6Ysyh8+1Fq6OHMJn4MOeZ4pRkJ45lAr6TFuEFtLgkMH12iXxexxChAclYOr/jGnCfnSslT
tf0B3UwK3K0//v3sc+WBIay+3DySDefLpF4SiYLqfySz8tpVIfudG3ZIFs5eNhTCzZTR7V/8IIgw
P2RiWO9e+WnymXnINo3p+wKx+bjapPZmAdvFoqsml1v38tINyz+0lkdgQxK98/L2v6DiGg/+l4n/
tYjrHfm3cBcWqb8k1hbY5lVvxEUGPeVQ+UwVzlskNjkCKL04GZlNKF3CIfAS3hf4D4LqutzJW+vE
IETlKkPu67tWqBRlnq3EJtv/guQWX5W2xgCckrIjTdcjkAxLduGvVXhfcIcNnHm9w7rIH7U5l0qw
aHLrf1MNi7GquE0XviMMZDOBVfWWk69pH2iLk+e0P9quQw3h87AnBOzC1ubmkyDahHHJo0GEtQ9b
JKSvpVU/Sed4RscTnXhZoZzjF27gqritnkZPXCPWaZQAlMseW1HiI3G8bZxBXPRGgvQ9Hr6EVQ8g
iQeMKDP6woG9BGEd0D2fkeruytY2JVbatFp7HhS2xJ+C5qVYENv5RJjNMkz+IN6mipFa0mNLdZC5
yAvBmKkfwNSCskhSkzpImQB0yxNP5RxAwLKQa7lX8Q5ohTohypgy62/J44i9537UsSoT12/wpZU0
NpuhE98Aa5piA9mygyL8GNH6PZUePXDRNC/V6esHr6uFLoZZYD6begznEnLFtm2fj/r+HABju0Eh
pQ0P42ktHHRxUUqsoe9fs6Cvc/deETeDyLrXXtPS5S2eSUKWTqgjMTbL+e6Yx3Mpah6vBdjFDF4X
4XALB2fJkr2Cky1gCNeXVElyhLA47Re1GENzTqYvMFgXDLgqhGlRBVM6TxsHvBze2CmlG2PeOgSf
MYfqrvLMQWPiX+K1U7CkRdtjadQ6VllJyA0ls8Wbg43GQkXYVL6eEAi8anKFMv+p5Tw2prKh2c0B
UrLXNElHCw6wiVc9ZbC6k+8RCF70MqoPf15pN7q2VIAv9MtCTQSOCHgVCJ0APMk3BoUfHKWdC+79
M58yD8SwhcJu4jdHaJKW3/t+5DQcjIDuaXWkNhp4jG8LzCwrjNUpBLyR01PUBoA8/AHUXxN/C6lF
1CQH20sqiDSYEVSXK+OhX4B7WcYfTbAy8q4BwgyQxKN5yT9gA3HyHXF71ntMX4QpqQBHO0hIHfto
4b+PGGfLQ6M1fpMF7jKIWq9hwBboG1L/hPpy7I0yIkjDOvts1q1kjDef9JzcF/WJAGfjI7isOrwb
xCwvLFQqNNYIgub/7yFisTe+d8ZAdK3dRX8UUdC16gNemstoPpTE6q6dbcD2oiBdNIADy/G4X/Dc
d6iDvboT6gSQH+tADGfXdEBOrraHGFTN5ChR60R15zD75C2GmACJnrD1PD6QCXdE4rkMCpLwmSMC
r6w/4dzonvox7Uxr7nOJtIHZmjUG/SlX2STvQf4FSaNPmY3iAsBKvwL7Zt68OO7vQIpzATwf5xP/
cVfAzKmtXgdYKyTGts1i5AQYGef3vSzDMM21/GKpFU44pjr8TlrM15JAlLAWPCLC05J2JRZf0o8x
760mz0ijnB98XIn2Vgd+OGd9kzZ0qf+APwf0u6shxRGdzBg67PFnAPVU0XYLbwaj4CnyVa6Y4M3x
bJDtKacWAGWTzVoEVvg20CZ5QPlWOCCnIqrizi+SLiFzmqoCUTOCCZU9w5v1BZ1R4lPtQwofUtDs
8qas+Fg0hH4kA6FwHGUbfpIZlNrb42zlBrA+fNOKbi4Wb84v1cJXg6zjt+CeFs6w8fDdrhEPcBss
tM1Q/szpUrqaCZBTb31rBJXUqKSBOV8bpsttTjs+UYDWl8Frt1PyGw8DB5orDdWeihJr4JSnu0Mh
+nZk4YI1Uk11/cHlDNDm29gTq6Q0ciYD4rzO5uvNNmdx8m+T4h7A9g5MT3f01Cb0Bdz3ngiykpKj
8WWYyGL9oK19O+vcnTlFvMATnmnqLhy9hJ43jvTN1PplhV+I7p1rVtRDe4OJeD+hAE/nrwUSUCWv
y8caPtidCxHHIHcef6fg9iiUhcYVdHSHbbu5RD87AYl23XkXj2CE9T7BNucQEmni7jnR2e+fvT0k
SrvghXimPRrWMZxAbZyveDRP+rjmwV6opqGt2NPkVG2owsDlzFZvOfbgiYKLM5U3aghRQOCalfL/
jkbT5VVqGWdB7oKIkE4Q4I3lYPoBT9oldZNvN00Dxmo5S9HFg3Rk/ZQBq5Vk9HUDklCK9/bv4Pa2
x1WqouMSEU1iN0fAkhMHoTesRNhAdxN0Kc1hSfLvoEwdnjFqf6jRm851x2dZXoytvUox6ptYExTO
fzHSgBpwjrqRfjDMDAzpOqkYlH4dWPUbRFrLdljWyjyXpyByqnUq7FS3y0j/smXCM9kzlTMe4W5M
1l7Wfq7qRgHlWGHdU8m03k/7wGKcO+4WcHRj8ADkay1EVE5QDhzB2x85Rv6BbMkCWclk6ebsZ8jv
XmSaIaLuAppkZuF47kxpHht1+xeTnA7C6tlQWbx4WRakBZjWfdnwUadWz9/TFoSM9MgtYVeTfMYh
+j8K0UxLP42eC+WUplVjdv5jUpkeA+Oih5+I+MQmTiDtd6SeAcS4z+11rTHVaOHSXMoxeN/axS9m
cd35sxgFYphXZqLvS7DPKkkCpIxPjZfIo8jdIQ5tKDd6wqk3BIeUv+NNw/JxcBluES/JwQ9vrtLz
sDWJx+zlQlJVpkHyKW9DJXj+c68OiWaB/IkPC2KLtIAIfmZhG90uUjnuqElsc83YLIthu+d9q0jM
UJnCEuNPYHA/5ReApxhTvhRyZDI7aSQompAmYwnnx4di65y7DN5rWx0DY7KJgtAkhqCLs52R+J41
59txfbmBqvuSpXvg0J4J5RcMOPneinYtbVrFEmjixQE9JCKMHStKkCtVTn1MZsimA7k6tx9QXcV5
761Ojp44Kky7WU3YY0w7tHGvmji4ejR6qaab9G+55rNKJn1E6JtynNTFLvg6rdHzcIO83JQZ4FPy
q7fitJ5t0vPqJfgCbLxWBEcUl8f07rqDTThVmUSKNcnIS3IF3ffX+vUGeLyP56UolkM+3rsAjhZI
/uK54R42J1/qUjNwgtYWoWM9lDt8bpfD7lR8nICPjlqrSoC9embnwOLq4osEXKCE/9GmpzXddaGZ
F/9wWEku+gtSbpiskZNCMkrBQo7cjW0Mi+LyPB3JdBk9WgGGKtRX8oD8uvEt7iEDqOUJf9OlXAG3
gnupfRXuiiXd9rAqG9zF4tahtjeT+7b21v6KshwN+vfLIhe6JrLRwAvYqyOIB/hj+uLaGMEvgmIz
+CYpH5ewJ4aQz/SXSeLZuNKYSKYzR1Dk+PGYl+Omok+7OuSburNlUGwvjVMzKqDNEI4H7koLsiwc
icRvfRUK7OGjEi2mmmvEme2ZwX2NzvOCdxGlxomoCBfyNggUxWHGnv/CiCF9IZo7G67+xk/L/m4Q
zJ3xLsD9lyVClmZvH/IUBHa4IoKEmVDOfzeCmlzSzxM39OHI1ukwTurjeJ0o7m38XocAdAVZw73H
/xTstOuOg/8aI9tfdvzGG4pOfreS6iNp8hh6STZx5dJ4Ti7g04J0MN5q+MoeFFnHgeZ1BfKjJFir
D8gr++o8l41f/KBhHjoBcqlYOWc22VfX6X96qB6DAKBGBC08XWA/yfUSsw2sSCoYiaJ0Yib5GKPN
7YmsgwbyFH2VaDNqzrWsnTi9pczKjtkC1RILHL1XS6Dpgu6nYgcP4Lpl4HI6MNCwe/hbovNDGj6T
hAPCDw1M7HFtj6kWo7nioHdaQU7HkPw9jaT2BbCq2x7M56aFzv31I25ZcUTksx4aabmcU0+AOyXh
pT1spKOZ6ytBFPOszGApqinIPbB+cWrFnaWkM9HIsgrsBnBNVqzvNb1J0RzDc5+WKU1VSmmF3IUw
X8njjUmvj0f8lFgQM1728QilnciUPXtXrZXtjVpaWnkmCIf6ivuMoL4X7NU6/3Hg49KHcXltxPmP
87rBtZ3X7p7LtYwJypL1w+5DHbINT71GiVlijmqNgUYPBwGUFmrJaFtQYWe1llEta9j5jYvXjubH
+HimlTovZ2Av7YIMgOd5KWuGIL6fkyQDzfN4BrDT8ZWGhZxuZ9pNb9mVt3IBpSStsPVVfzA9TA6K
F7iEEjLZrTye3HiZh4p3aRXl65pQn9JJFwHpTeQwdD9NjXjNa/cgvdBCd2ZfbM1LrAa8THY5ja69
pjWjRgdixMyG3pcEmu3lBYELftul6FcG9riE9DhET296hXt71k9FA+XUO2bZPlmw367xHM/xpArW
TqP5PGhWiEDW3baDHcDjLJoyokTHg/OxpxLH4yMyG+6LvMPbnrHOD8PL6iPWNg08N9idiqS1PFDs
dcEQxeepql4lEsRmVwb4Yqvb1091rkRBSrLriXGiC/tFVg9B+H3TStsnvWokCrc503Ii9Lg8C8yr
i2vRQ7Txtzb8KgCChhiQ5yxLxDuphLbUXhX1zJIUGlXyTFwMotO+5njqjHHBVFYNGsMuphFgUkpu
XnToZRc6nEVWPQJvTtPCL7o3ImK/XHBlCfU0mHP8Ov5Bx4ELzPz5XP8niD9n1Fec7tJlXKYNpemi
5OyAa3Ms8f0ZnPhK8Mxs9DXbzd/SZK00MLNYCdbyQphhET9dSnjAGROrYa6EVlfVUsIvg8+DsOl1
SVmoZ4b7QjZnihaNENfiYjhSVp+whhccwg/LJndMGxLsZ1jr+jNyY9Ew6upLcdM5VTkOsLGx9+kp
k8XoxOLsqjYPuIZ05o8C91fSEfQODoxikdbqRBMWa0hcuMHU3I9LPCx5pky7N5dcmUBbYGX2b8Wn
rPAOxOez4cpLF7OxiE851MCzAChp/ZsGeOnHYUQMPYKJE1vKUYBEMErHi/flnen0tKaSWsnFkrtv
628IXZDjQrQluRr1LGzv29VpD9u7EmjFxKVJ6LdimYcPC2ggdMMeTlaKoO0l58glpwm2WiCQhBf3
mYvGTAxh/Jygtr2AK+HBO1Kj4O2FRteGL1O8Lm1HyDncCcC4IhLJVMD6fbQSv+Juut9DTtBJAqb/
CSWZYEGaBrVfj5pqdA2CGREda0k2w9UylY7NPtGNo9M3ncaDQOGUo4pmV5htsm7X/UXTjdB1fOpy
5ESSypRwkpGCKH9dk/urAydb4TqwQf8rEwVZb1RNuFm6BhT7TjO1tzJ5UL3WMsAOrAHbTRHrs0mp
IY/R7Y2oDJIIoukEU3XEMB6ibDWguLGJLzrBE/FszJ1DbYvYJU/IhClZi3ufUZOJQXVVGjYbHit6
Cc1rPHjW8uFclwbL5N3Tmod5YG0/r5hbxNYeWwBxjjenX5WE3wJ9Ts7mrIZBT/Ezv6W6WuUvCvD4
Q0YyGET5TNgOzvjI6ptf4DmXBtpPppUY2jH6OXd/gsTb5WThTUs0mf7Lx9NK7qDhfl/E2MqUfBwk
bFLD+UBIbslAr3Ja5l2RuIwVVj8njp01RJw6prUYedfmtucO78HMlr8Lx/RrNYRLDOPv6ZM40xzc
M1VDhbudr/l86Jw0/hpajiyXH2P3+8WBNi9qGPuotQ3GLdcbRU5nQg47H4w1xiC3B9p6ibvFoDT0
tph2gbE1UcFIUt5ZVI/+m6TcJe2mhjrEQk7Aa50iPPUeFPdtwCf2+huwyezVNdNzrXY9KX8pgvhV
Z4bel1X0xKb1ePvI9+KBFT2j2d9RrpDXJ9ue9Ynlwvc4Mizth5IK5sKPTaMQamRZNihkZ0z0KPOA
DXkuclGcGVLDoo1C2mFUABcq8NhIvDrWTlHKWetudJOFlVujOULdmun4/SRJ0vzsXIECunoxAwqW
mZryaFggMoJs3sSKbfTu2bvPQB33XNUz5xo2N0rgsawDxnPCnoNYlVJvJSvekfQi175LqyQMm0QO
tsWxoLCt2IZyGfBPyZNxi61eElMrxb0dJtmXD1XzDQ/70i1ptwPKD36oh08ZcHbbLlNL/rILkgME
QLaLMUAFbr5Ha9tp5JQE9yE/P0tnNxbAx9/sbLGU6SWCL/dpwSW0/9cqDw8UdY1Uo38hl8c+4rTp
SHPpB0LqSU3KurTQ7hJ4idGO/uDWHW3RcDpG4L6yEaS4yLH7t/fr1DpXydt6oyXredi84V6YiJqD
V816HpjVfudA1PeDtvFbX/qhWRd7BXvbjLvY7E5dTv8mNGLZzqxjjQ/XiJ7vbkZzz+ufpruODEUk
bZ02u1L4tTFvrg2dE0r1G/wL+ABYtpGug/VBcjCDEWyDbRJk85L1XfbHbzx8pRQ9/jUvwkE+Awce
halQvsVl8oTX5XuKj4vnM/QO9YIuvoy98qC94jnLEjDacHcuYlYYNCatVUvfTgEEjwKz4tMaxaOv
5/7RlfjVc6TWngaEIOnouMwq++ymriycdkosCCxRpjxcoXpPTwInDspD39cuv5t3J6D1SAWMQhD+
gCeZKjnFm6iP4wiUQr94U9DtWZ0j2kD0174/bhSneNi8tfPKwvKNUTm2+uuKdimWG9TlOB+TfAaB
oJ7wkCM1rt5WspHdZdoFqpk9vnotwPLdUEwipq8bhWfcVF/rNMz31IgYig4GVLggbVcIY0R0r+l9
tZF3rfBw036cl/zlnUR7SYwOV9A+mh8D2fZdMyke5HQTEIArFeRYUrj8aEWuO4YAspF0C5oOu5qG
zNiE0iA9BAFlrtqgtUUrnPJ12jHS6e2gqaaK9ZTrOi3WJElqZBnCb1E3+LCYka0xcilAl5vhDxSC
c5poYdKRQDTuCa9FnyNGxjUkMx0Fta4dIbVLogNGtj7/RQjjOuHqtnKsKmil2lRX8SjgOcf09TJy
gdVEIyviaYH7kiahFqWA10I3dHsEWN8QO1w5xTNBjCt5dvup+KqdUQOcB1W6EkjpEwNd9ElZL09Y
XqMWw3PI18yWDE2XV6j0MKAzWYynveNVtdznBHjIkhfZIAMJ1xKOGKRV/JwZzrNltye6MHwR6U9B
V5uue6capfU28z9LcK1/ugr7MddGyH9wKAnzO6Aj+zlGIeiPvXB7vNNtREFmcMAAYjNT6fzSnJTO
9O7OLr9L0VcO5G7OpVvyAeOEkyw79bZDGlGPawZX6eO+eymPlcKzaX+JgEWAhrD9RUmF+VjXJTEz
3ljB+ekOE0IL/s061oNMy2xel7OX+LEGTnDnhcxJNlqNFUmKI7eePmwkOZX1RTNq+TVNXoyBHVlG
KapLAQahP935GA23AY5ZZbvZcMKVRS21gUpjbfDdYFOHFDMgY6xBUCQTSIQ6tSxf0nPORlsoGw2g
f8bmvJl4d8HV+BWdNEqTcNreijHErWiZI0i4Lf4nzcfPjrtYg4xFjzsO3ekx2rqyi8NDxU8QJMPI
nBFIvdUcLQZsyohZFpHPWp4gXDbwOXoXTccsuLuL4n3StssiYgc5VYlql5VAyE7JZpZu4OxH8T8G
rNuTtDPStKDqUtN1hvyBn4HggM/iuSSwS55j674NOd40pmZFLiuxvKmKbcAGiSLLjRB+mDgOygV8
SivAd8Q5diZQOf7h075FF8Y7ualpwE6a0PDv/l/nAdRSwy6JVDTPz/SCUrkBkW/Q5aFdXZTZCq+t
5fjWSDDJwt+dtPtbVoq62333beuM18oY5HZ1oSLmbSxCbm9ckLMJtwVXma23SGwe8koNjVylXptf
1yND9V5un15rK966n2HHMS09QNTSFq11LT5FUDas/J7lV/kGTT5PxnMyG3mM2iXyvOUCRIdhZ5Ui
FXsuV11eKB8XmK6HLPWA18+BjVEL6kdhrkRN1gkLMgx+isnhN1EA/a3Vn5bZBII8X3/B3Fv9pRyc
jLLStyNrRMGWn/TgTfq00ZI/8treQRTxSCZ9Wp/z8t4jsVNaibjRDarospRHmmJglC3PI/31rnJa
UKsDXDI5x6+GesXE+G3NmTdZG7aTZBrziHG00uE60s0xsexUjCNx0bmTDWZHq6WmCn8Yc1L2s7Z1
J+gkjWXEokFMWsMSSjrhq+grtZ7exMOjkXRSoaYUFBfWUvpBwNF4gZFgixfEP33ZZaXWB6yugQNl
itFcM8vLh8E5JngWXSPCtEUvy81YsFHz9jfoX8i3VPbiYwMubWUto+9n0dugv8L2m9U38pf/1RMs
qkdmsJXo4novZ6pov9ULT85/BgUSfO66qamHo0D1Td/4kaZy8jABzitSLc00+A95Hvw9mEFgaleP
ZVLGZW4nvg8LYQdQfss3A8D6flDAOaG9Uzdmgx4k21ibxTn1tC9Xy4lNkUDJnVXaaPbuj2azOL8W
p9vFeM1SpTMcN0EUbrGqaZg/1JKvbKxQth7NzxPLREoZA5XP4c/F2XlhLnikSP7Li7BYDa5dlnl4
SdB+tekGQ+OVCLr46MV5hm63zoqosGyCrb4DYjZQy8UQWWb2Bdg3e3OS8gJBLTComRGl4dOmmEP6
WydrnmDMRHkPTBeTBt+Yy4JC+a/sD/CFIA74woxiCpHBKx6GM+SMc+71/4p3En/xUOsojFCreUte
7xFAO5F0i/XYod8/G0nGFLRxx4eta7g+wOh85Y9KuMbG77Vwyjxvn+MF2Vtd+dSiacp/BuxIKCfH
KcLcOzWfPmHDKV0tAIa88TtnkRJN8ReJoOcILvJbOSDvfASq7V0NJPIbO7BUgX3wr5i+kqM53Blw
8PvPQv46qCpy5UmqeQFvi2HCzME/Ugq9TIbdjyuvR4P7n7sdaH4naEJpZaDCIJBtUNP1M9A6wKn7
sEFmLU0lZ2c5FGzfmAVYj2+t8sAdz7oEVsSAfUAFhBZHDuYDvUKGGW2etxUcSAhZg9YaKnjT+XD3
Y5o6Iffeay8KYZbrGpjlahfXdtSg5NnZr06geXhnngF+l5RCtDoxjC9ON69lkrj9pLq+xlQ/6mjq
zC38kVQznArjQ9oXlC/fwXncpz/Ga2+n97J0q1Cy22kyhIRrXMcrv2O0QIE4ksUir9oLQ16WD4VF
uOQwaF1zdmJeClBHX6CD0VSs/PqHz1DuRaRwWAlpDoofgZ20hMKKXzNlGeshm4KsQ1XqwzE1k47a
WzAsLBwqKhxvL1SbrtI1Upg967N5u8vA69uHKNoRMsB6ntjckExlCcD+J7LwDX4NfoTcnI6xlo13
NihfiVMdpMVKGKvfIHCMbXoBHz68EEAR0E+uog+i+cyNsrTCcKNyFs9U9WL1TT9FkPCxzhwlbzLJ
3964ElfFzYSo1QLQDv8y3umcJezvf+s7Z+a3qjObK6DDMh5hy/o1qJ+Gi9SvHwJj6uNxBQ0Iuz9C
DJsrBrL3Qj2y0pyYszeyedTyaBTcr3P9lolcAJdM04DJNvKsi8N9Bac2ZcklKIi0T7v/cMKoXYsR
JTzbH6eZgNejqSf1HwLRb7/1zLbgexCEbgyYVy5zwXAIP5hrSjei90drI+taceF36O/jW079IaRC
5AIQqWcVj/rSf1Kt24sfQDlIDw+FGdQ5xcUkoX/Jx7M5acH0qxS2JBkHOuPkHeGO1Z8/o+vpHZxa
7ADU+/ESNmjHh1cP9oTvb0lqiiTSGDUFTTNzuGaK8ElLdK48jm1qABH7P8EN1v4L8O123iPOisPa
5x5UwSlEfyVVimZ0YifQwg48j1EXoF5LLg7zGpGzoKy7fUWN/t7FPPpJ2y97p8Xnl7JhK2a+b1Bc
hPI1mfS14awou5v0svwnxkRqABO9BYEbbhfOPFPw67+F6CfQTHst606UAvMADxC35zoDuBNqivug
By/N02oQSqwiZXb5nsCmWRExmFETvNEQeKHb/EvrjJippI09+sF0BbPYVGuIrmugZ1Gv56SECEfQ
fh451VC/NlHdQUgkIit1/wTryMVkD05kS1pPeSkgvxlwYuzoGz5ImIzTup6vKJpW6GkDYZGwk3at
B9QN8PrqSdspr6y/AEEdFtpnPozJ81EOs93l0g6prWRTWkkO4Tuyx4C1aRTpNvYcBgxhbQOPwjFj
e5T1LfPCvt1SH8RhUNRwqzT0iCKQVVziHHS1axF6MnM39p1FJsUnNemKe2K816/eO3BVuTAgAWXp
zlNmYUsuZ/G3ywdx5y1kyK5YWM/q8g6gDNTznrfKRddC4re5uOfzsnmEoZDLOM1Fr8MkniBpwQg5
n/U9TLC27rpSB36NefArIlkfe1RHOma5r7KeNhYKw0R6mW0ATjvimT2ZzLxZyADUb84/dG+0rC0/
DkPdfA04qfMTuLaOMF9jvrL12u3G4bWSmerJ0kJh2aE2GgzNnY9NT0bgNeDESPbBbWpp+O9KsKUL
hbBRuBB4RiIpghx9leN2UQwZKPGDs92it2NTSGRe0YIZ3EkZYUu7bThIRcwukoZ3tl/6XBRmQ8F1
eOdFG+naSXkxHMVVfUVqlsdXzLOwhbMx7d1++uNYtefg5Bw7pHziBpa/GTsaMqiqzVx0XKYLV6Ln
zsh3MvQj1NoQp7Nn6sxWg6vO7Wn0qO0FkyLr7c/35LlKkIqE5Kk2Vr/ng+5Mkj4M4F2z1IlZV609
k+L5axSQf6usxz99W7SMhEr/YktExjnWcy+40KC8NTy2yvK0ieZfglivCE9r71vnzNr5KAFM4mo4
oTMQzkKa98Jmqv/D+H8v0dHYG5oqJfr8I7tkislZReu0Mi48A1lO3SkLrxm7lzx2xSL6tKZg3T+/
mMmdAUIggp0rOJ8cBgTy1BlLREqWQJbSyhT6CRhzpI/RJ0nCmh5TiyFDJxBfUsPYGHg1SmCKOJoL
T3HpPmiPJFvf2GeyTLTlG2ymzw8/PRqFPwTh5EAZImcJxGdwhO4y+5QjO9S5r1YlFfKdrR3j6wbH
MUFeB9QwV+P9qc/hMPwvtbl0YqCczx5Zj/wq7fLMOo69aDl8SvVXXmDd3Q2autHvoUqmbrrq8iW9
PkXlrrw8Zomrisk+HvguPp4QHRvcJmWq3aIECCDPkZkVXQB47gBMsm7KDgvcCoSaGqqYbDqqrlkz
yD8KVvj+RrUKV1cOxJ3yCcHJul2jsYIqthwAoDctxElQSolpJ3xHM9Ieb4+3BwWrs1q3kx/RdBiF
cx5gT6PuzQOzdCwYpwiGl5zqhbZlDbc8j4VD1hs+qBSp8Es5HgdzduR+zrM7NRGq57MOWpeEfxaN
VzFjjkI+O3sfmwMtd+Gs6h5j0iJsiVMRKL88fZ+iJLVrrVdhM/8O9RaKMRXWvNImPtzLwVFLbhBv
UFn9cBEccY8n9TN0Xx3dpBRaHYvdLoFc5KMk9cPmLTkhbaqv0iOY0QCraT07+5Q0gd6J6Z/kRsR/
RNCtd98WSBS7LYbPgQQm8RFeoVgFWo9+IvvtRxyewV4j/6tOct2AQeC+2G45HDUw3KXaQfOJQBi/
m/IjM01QW7QZyj52dXJFlgmi9qjW5NPI18ZQjTO4esVHZjcX3xnFrlFCSyWkCA5/56ChWbPwp+YD
aWIGTNhX2XMmL8SfK/5+JHMLY5/wqDWUSZnc3dxhQVf4Y9fFWmEI7HOO/nX+925axHoNx3zzxRr3
lBiY77qwIrSGCr2WhwybcsjEsbEwePaszGoRis4OCOmMBR29HH0qDP2FqENdOBTiK308vvDpwZ1B
sEvXt2NPMXq5zPieryxihWkSYP1sUFrITt11HIxl6HDd7m+A7h3MGDgDiG5oan2/4Rf0/NE5Nd3d
CjhwrJQevMyizr359YQvZm0e4M1mRpvaGcG0fasmrEDXNjGvM33GNdtivdZpzfJp5j8E/5eS2KoS
nQdiH16w3qCMBzMDgtzB2fKolDIwud4ZneAP27wtJUj8ZGisXW0sCJn0Mb1LUCueDdP40iJ/E5gl
re9QscabRHxTfVSaN3bYJky8buQnKhWDEiSF3yzMZDNWxwMKLv5+bqgQ6CJu9hmlj5bm7s2omybm
awZZ2NWYpwjccEwuiAWYx+QyZOroTRPI63CI1FvSmLR4OJbBrOwNupcwhwORL8oB/7TFUWIA97oB
pVxvudDKCWpXOdU3dmPrYQCgb7DhYnKUxUsskH5TYVcVoblBM+FyKmMXAzJMzoavFQPon8BJGlGf
fxLb+JHjRr/Xl8R8af97b7IL/iKEj8Y/fmUpzaoAqUi8d4tH29DIs1msl/fE0oR7omt56gr+v0k+
7M0g2CtzLpHY3n+Y4gbS21d+CKTToIzvmuZq9bMTYNbkcMSfvBiDSUM9cA2b6zWTEF7BEvhhYSE9
BXpEP9Dg4EGBorXuYd6pylZwiXZcRWn2ZbJcdLLhSUv0WZFf5UE15E+Mi4+3Kyo6ObaARXOWGTy3
/U8JDdEOTUeA8IWvpnHk3F8i6gxU4YetTdmUM2W7EKm0VOgSVGTr2H4Lz+zqAO/nfPEEjYQhZS83
UEmo8h+XQgkwkZ+EENxLOYkVFH40/z6KLGUQytgHLVusNisAZEFWOQi8lbS9nnvfgxgGD26hEcgf
LY3NifNJD5mImRY6G53Q8VtdyQA/8vxDpB0PlIQXEUxf0d1UgBPVaGjYnykbuNaUmFXEuctrFrRj
21VRKlOh0oHcstEchD9BQ0t+mZ4qR/1pQ/+FELG9yWP3SZPMEo12j+MqWmU/r61fE/R3T0ysw2tt
0dy5bq+d+2Dm89gj/btU8byblkkdnE4DyEuAdgsLkC89HvAmoy9qCGeyx+dfAUKdWTp3Ypz5yB2I
1gQVcJTOzanIAy7XdBN8xzLN68IMK2BYAYkRW2NLF2qymyU1avTFbzhRje9EUSu1S034KVtAtWXl
WMXzuyinMusVw8XdzX0cyct+bu4iLo8B3H3eyRyPCRnw8d8ZCogUy4WsoC2eOCbrEYFt9HY/l3nM
artpYbS32zIForPphWzadccltY18yu1dq9KzPJ7Jtd1+69za7wwFSalJVOaOBF0sxQ/7ZF4y+1Ny
iLfmJg3j033SAqCAbXuhrA9fwBf1sGC6AkTtt9Kw+x+92nkj1Gfpqf3D2A0YcbLxzPU/X74b7aZ4
euOM1cZLAvtis0Z1/0dMzFzDY4acR5gV/KTmg+/ioBDyagJvOvYE1+sSQgBmCbqdeqWJo/dd2BYs
GLDOKU+n7MnfxySWVqY69wgHFAXRN3Th93MPnrd31wGCUplNhV/rFHnWvWGsjhsPvOYE9AzgSY7d
tuSaxLLWTkNajzHZP5riPVf74rwOhcNi0u0gwXvkc83Kb8H/EWHxJM5rGrQlcwDb29TunNlQKI7A
LCBlwi4Yffk/+TUE+JxdshDOAzSGKJ79qXfrJlpdYnByM9HVB5k9WuARW2LTCYUWRp/ZO3hlZoC3
/5sCTBdMh73KbG64agpGhscTjD/Qem3I+9+Qy5G0MG+SkiZHJdFMrgrBGv6+Pm0fASptip1W6Qcz
3pH+mKofe6BYeKROX1V0KJSllrAgU3RnF6jgIDJP0/GTvw02XvESSY6qVWQgoJqx1NoVrcJYJN3k
WIBV/7nRLejhLnC3iQ3BEmLCSCM3upq4MvPGWfu57cGWmm6xS1zwX/pkRwRp88cL+0x0AhQrBtkb
1JhPMLkEwH16cSbVoPJHKHb/FxgSZ5JqKwaYoXWYGii97MgnKtdhTuTbBnf87E9LE3Qx2U51o4m8
yrW8WDQtYoh+OILaWmtgjp7tJVU+/9vDKA5haWVtAh0JC5tzvaPQiQXZKpBBJFw3uKxUJsCL9K8M
fsghJtWY7lW6kNCmLT10Jxet5+koA68RMP1J4f1op5yFjo3FKA2HLlRvyaajXjJKhnTECQXD7eao
2yG6MXN1/un2GBWDOi+SbSs+jy1jPOrEgCWbvs1uJdf20jSQ/VY6KZA7wfp3O8XTyKoQhJ39aYBY
I7EatVCDn4FWMCutchSVzwol5htDJ456D3Zc2HqsL31nfp2BKgfPQrKtHnxsiphQ1cF17iJGTmOO
1G4nO0SdV7BbtSEBQof5rZj40oqTbeVL2VZDh4bkkmw/o4EfZK9engZwaAZs9xQ40i9D6GDZih/c
cMHk410nbi3ZET8p4OszuMmw6Akpuyf1Gw65aRM3fLiWACrKDKlQlP/24o1hS4holE6xk5fTR3lK
9nJxDeYid6Ir/J2USSmMR/weZ5p/XfjPG2Uuv6PRQLpDiWZgaLWEdAetEFHq3rQ8m/01ttpDCCeD
hqzJNG1OLNqo2zkyHnJY+fiw4lX4dVZKmFqeB36KotjamjzvDCPWqteIF+T0AgoeuJfboSKSauCj
qb5smnW2vS1bcyMPeDjqVetvuES4ut5aLoLVLJvupFGGRFZWQGqsDHnfrnUxP1ITLv4Vf64kjaG3
iwo57zV2oxb36KZ4CxYL+sLT2aYXqf/k+mj2QCCEusNb6CJrmuvgyrFDevPmKjCJCrcDc7x00tqb
0gixlhpWNPOThEFSOpaTWpZn48B5KPIr+gr6uHMxXTRo0fa/n1zSfEQ0dFHU7371vkKzagB1+UDL
8DhfO8Ch+fMvCh9iXqwWrhFYOpDAtVMs/Zg53aOZeRmHTKVK1ixPkmq4YGapS8O/moyxUwnnjsqi
vos6SKwtzEwjApu4EmT9T340zTNwelmEJHfTSAZxGc9uXWl/q+bl/XFbdOEVTntgwxJVgm5oRoro
S/PgiyE5/IZOiS6fXnHkplLNV/O8dDXKy/iRvCfkZD3PupKEs4ZoxZ6cSbQjNYZDMaGeiM4ui+DJ
IHjGabNX8HsQ+WtJiIupCcAv1gPStwOuRPYjzUNAFpDYnIxJajxzFXXzF32gYBEGQ4kduN6rUpey
OK1lLnHNCDh7grrF9J7cgx+BGtX2H2Rpzzf122tEWjqFPA29bz5eF+aqzC3owMMEYAlbJjgr6ZBP
aXhlGZxMNSX8x4mdeGoQu7tUko8K8qVZkwNhtltJcQpQPRtepBMnet5+JHds9Ll2Zfqkq5noVqop
VHQwRgfYuALEv80ahJtUKsgpkTaofNoJbX2VZIaPMWHyXRW214K/4OTVd0eIWa0GXPbbP938dEt0
2/mJSZsfwMjJy5AhcAmxB2gNwqjErbSPGoR8/7YdDH/92nrSlU2w4fbqXWw80/2JcznKzZTUm8dS
jVVKOBy46GjJC6zB8ATHZYihOg7Fmjza6NyriTC/009Te3meA5cT6Gz1cNv3BPdOjg67fSqhTca9
PE7lXggPlCH6roHsq6fHAX4s9HxyuOO98KmfR18m7zCjEFduxuPnz0FoC2Non4wKM50JzaRvOcD1
YBnDrVD0STlv0l9oBjGyeDkyvwi38ArJJcfAjS1m7RI5CmP7MVTJnQW2vQkC0vzjj9S53x/jEHZ4
3wyoj0jgys5t1mwPwNxrKY0qc5ZIK4zJWvrm+DxIi7PRrPA4cAOPVmEA2BqgM4l+7/RrwKkiJRwM
wJL6CeDO8RePwYj3xun27LSisnCOW71ZbUuPha5vAlwoB6ezyGsGNPjOm6T/70EWDhNwy8jkkrre
vw8KuWaGgQvKdQm/FFhCyh8/rgwS4IaS4CB1RCC/E9Wvf/lpfcQXcgLiF9yDNQmkv1LuRaHEAgNu
sqYnFxQIrhExvfKhlZpCnzVMLrE+hF87BX/F1bUqWV3LE9ZraF2J5aJNWB4ksfUrcBjrcsmMh6LC
EIpmjQ3eVXf5OnTxNdtoBbrRTYXe6qWZoK+NIc1JMplxlXRwAEON2hi78bEO9k2LPyrIW7NSsGeP
XZEmGgqn0KG7STF6qxEi6l+VGxJuQD80GJLgkkMUG/4O6n0QD9Gt03NJ0JYJcFzVBxTuouk3fQFt
dKIMNcL5DAfO5jNItnYbywZZLbN3169GeQnUJlmPuxHYp7ABk2C6qYztL6dtgftHh+dZuZdqN+zK
cC9GJYUOgHY3VseGWyKcqVolRtusoahrJEsLknOfbfGTa3QshFLxlMt6rkeLTouDXPVhvklqZYE9
gRoAjyvcpkxlLsecO7oNoY0mLBF0cAoOZ/LYdRdOfbyX0s/BZpt7Qj8n37BILZf3r0chrcoswg6K
Z9lnpkBUWLgRq6ktWEbXD4CUCrlBy33Cg+yUdOqAFWqVvTz4QjX8D2fNJUMzvTBDYUqUHUniJMyK
8Wp0BQadbYg9gHV/ORm1OBopYRQAYlPUekUnpEPChLrJnTX0u6mbOa4C/3Mjsk9ZK95dcOzsZzSB
gLDRX6vI3+PJP/ocRjj2ALFkKUJKRRCitGj1s6sEX61mZKZ8y8Jcfd0Wh+6wu3EDGdyVVMzd7/tP
ETNZEg1Hn+DOq/IVVFWIRWIj0Th3LlP/q+Ai+PgNuC7OBr7VYfKu2vbzotFGf1RxpYivIqtknFUx
7/dUcJOxskN7u1ZPFEAaSeOSU+NL0puotKVyac+/pCngJIIXV1eM3NMcYtrH4wnuIFhfcAh5doVO
6/w4ZXkSqOGp83DkI44M+74vI7DJzXW5g+7y/n+VGobRBgjKVYW2AgwQj6Qp4tXJ2G09uwOzPTC/
u8iKMxv387Iz2xl3X7Jh5ck1lzIJ7f0ClsNVpx0UNqoB9t50cC878d6Y7GloBvFKF6pbQI/xpY1a
i9C6/tn8siVSHnwKuldTdEPlrqhiXXCCvJhiEd4QnCNdTiMPminjrjRABNL3WbP037yeFtSumxXC
BQO7B/PNufAE0aBPzYMahBGXZvr17q/qs+voRMsOmNS5FevS6jse/QknrpHtvO+0FDlRKAYRgmIj
dzKulgrLCIEdj+JGHeGh8Ouy7RulamqeQB5X/HG7rdOv7O32j40uPUME/YRegnTV7LRhjXUKya16
3YUK3pb6ksJKlwWkpIlOekxaaMVCIALevhrlKmEODVXqFQBJEx+avGLpXlrX20HUSo2O88xTFDBg
lj+i31pUaNGJdQwc1L8qNNv+yVU2caXunLSztxh7kBf67VjnR+shcIMjIz1kqOMzgV5Tl2y49wVV
LpKSxjd/RCAmtV1+6hHYHTiGq/YIyQwVlRTzJKIJBLyabw58lPOE9JD/WkXoqYCV5GUkS5amrbp1
EkLBks2FJAQYwRPYA4u2HKKXilPMg1Y/5C7kUmZZz3EVeIhxsw/NcTu3RHpdryJ+kNU3/hOrfa/A
ZmImtvScUv4YDOn6Qk6xhcFAn6E92AFol7k/kHBfIrjELPUmS5VJcBh4PtcKcTOvxiQTob+c8bsb
MGJ6HbrgPmTLrUvXzKzlt5u/vfkBK5gLPvwZ9VsQT7XwSnlj/bEmOwXI5rpD+A+d3PTFKoimf8tb
wzOgYlwEhFSb/vj96QYCpzjohHcoo99R3A0NP7CZsmdO6A0Rv1wgfEQtCH/seYQdBdB2+yDK2GTp
rGbCeaeDFSmigrrsvYU3ZrzLFjtWXFzA8q07xJ9l4gRn0PRvqur+xvwdYFqXpqwfQAINYUcyH6pO
Y5MERhXYqn0KSjQxN5ZfasVuuumSqPVEfEmIljg0Lqj4QfQOBDz/nD6eAyEQxBLtoU9h8ifDjAL7
sXFZuVnzJdGNyPEQE82NwQweilK0OYmvBAAZv2WOu2nYo52DaXF/WUY6/VZtlECuQ/d8EH8Ko/gm
l+n5xZcBKhCO59TWAtUI+FXvYPyTy9MgNTIobIarmkOiIDiQR3kLAcCcN/mGEs9MM3ZDtgnzS50+
MCEpKX5d7UNoKEyO4BvG5eKcC/P0Z/WkHtfjFngLA/W+xmMTT+5VHLeIE4Bf3dyvbqNzTNNtaJS4
wC2q7T4eBGSDtFY1bPXVWh8yBgoZLydsHHTVJFFQKB8/c5mZfnNSU7M/wmDw+vNabsBQ208IXf/b
35zepbOEHl1aiOCSpxCxk8Mjc5EqAO5AVz46gZjnNj11lP8YaCl/iy2iPDExZQNovwBGcbprXnr+
l/MVA3uuYzB8J/lAPB/frZkgH+XmVYs3kiB+RvjL36oZaGl1D4vikZ6CRUxOMqUUOMNFU5tKa+cB
doppN0IEw4fuQfJa/+TQBNk++r2QusuRwCGLaoCSaXXdyNuGFO4JqFxCG/YlAC876Fdhegm2WlxU
t3ItumuvyjawVKmeGEY68YOyOJ/e1GzvJmAPdlz49lH3wihY6bwEXHZEvfUfZMyZSAwM1ZP2+XES
hfC+9b/W9w34PciH2tmDMAVQNGYI8fvASIQW+tUrwSeOux2gtPkoVP1X1cKotjaNGDgr6fKqOsEx
XXCsZbq6QN8iMS3+pEr4URvpQOWrAhwaIGt8/RKr5OF/c9sYVJ/lvBSKIZkauWnFhsSdH9J/rYR2
6qtnxONzPo6qm0KQOZZD4jkQJbodJLKc/c9x2PSmH+YHeNCQzgT2lDbYKCI1x8z+ObZUz5Fj9beA
GPbOsoAWNgsi9ooHT1LZmtf2v06/UCAw7vJKo0WZkwz57CFQmJG4m92yHF2BNRn4aysH+dzXp8dq
lw1O3k07LBn0ryHmMnR77FTiucf6PLssAVpZksuKKPt+D6hw2HgoaXrMR2Ir/NpwladMttp8fkjS
I56/JmgYvwKNuhV7OuS0uLKSnPLli+8g0s3bGAu2yTZDj0nOjI+VCJKHCUHYkkg6Nx2G9b+1IKMM
W3JRN4j8hctMd9M9QejMyOnIsrfqfS/Vl6rhlmj7MeD+jQtMA76VIduhBtOW1MiYQyi+Z03s/cyH
KU8egMGhWLjzUfsJHC8YOsj9qrvW3f1o5q9+nS730fNBLEbLghkbS6+/ontk73+YGsbJUKEc56kx
nUX2H2sDNb7frJucNRJqY02E1vTjzLDaeXoK30BxjNdom9nZwXQXdk0ELKmQRRIvybmMixA+OkUR
QsW9KqTacCfXnCjpg212Dbm4GdTBVaR3+NKJjObieiBmzzRfkYu6BHJeurSAneT5x7CktLbTJ1Yn
zQFTk/sWiByYTQkGgypomY2WR6SLnOrYIn2H31Upp5ulwQT6TNK7GHSZAzhqnmSeEh26ufv3pTqz
tDsRvU7U4P6Gj234RE1UjdHm3qFc53GeyQKseEQNCwgvy5snjAwWl2gTRbD8ueuHqK426NIjkPmE
7Xnd4moTxjxeEtmkiqlmrNdksYORYbUatZMnRF2nz+jV2+qJHTgBFaimMLLwr2vqMUYJ3QozBeBW
I3IW7r8/EMadOiyG1a83qfy0qT8ISL50GWLUYNK2XgewocAQ1sfP8fFNfqzDeFPPSkLXDytdUH7h
dBfuvfU5AM80eNWtli+bW+Y/ghqz7z68j6nU7hBxPNUbsV7kirBOnzfs1QvgiEk5Gu48e3GloI20
FTVH9qPcCp9FGCg1m2yRv/9BVKfiowPgA4z91vqZ2IO+0aKz553to09b1Wo/W1hBsHjdIa2TbM6p
u83wB8/NTKwgJsXbP41b83scIwoPsMPRP7EZwEuEZe3g5aHhQpoSKV0uU5wmqdBM+IRWh6wC4nkF
Q5gTKyKMZooec4hGU7jfuUylKXximfBvitRcT/xbxQyzKNw9s/yppjNVrMr5COGI2Bm/VRCbuyGF
EF9BkJBRyVSCvyCZKCPqvLuII/bEjwGlz32F+T+a1eOw2KPi4LVCDQOBLw/aG4yxYge3rfGa1Qrg
Qs939E/5mZ2+2GlonQyAOtZ8p/njykYgEx8vM5uWnz6ycIUtUF+3e35SDtNuROYYTKRki6m0FI5a
KwfozU44YirmjtsicYbib+0WPXI+DWbGNR1o01OrFuahLwPBtnjQLU/SokWVoPr72aFyeYGr8NuU
xjEO6J5WA5OZxZIEPl9w5TK7JyYqr4nmPKz/cMl4EIrlfZSxVCFNtPBn57REHt7LS66Fk8nI0bZ0
ZUU2Dn3R9OzqTWn1ZGSWY1xa+2iqu4quTWOIg78jUvxjAHsR/71674hSl/239eOH1adQgZL29OB4
VoBDH25ZyjByI51QvZ/TDTaGkrDbXNzriVgy1Tru8jZCQY8MrSvVuRGuE8kXDUnOXTK9sM9blIGH
1K1dUIWmJcFUjWQWOd9bdF5v7rNHdFWhU6qtq/zKXmMZJjcB4+2PYifr2q7tSnHx11MtOzoVDMXq
dDm5Ga+5Jt0Nk7IMjPmsh4sLBWnWzX94F1xwsv6afbZR9kwTw41McY5yqC4vYu7v0/HDfTRwBnAA
d/XtoADJWFnX7FUVRGhq6xZLYshjb8+WQXc0KZzPDK3K2vXJI39GU4NIWDSDCo5wyraR4DOpikJD
KiiOlYoqUBib/T2RV6DxHLLwCCJJSJ6REF027abCAoc3vyODCPYU77XJAYyN5tKW55vk4/Z5BZJl
Dgrsh/nNAAZrpF5nk1rnoFnuO6S0h8XbdR3N5HlbWIcLr72SZd3TBoMqMZYUu4KLlEcVJC0ZMJ1n
HidRUo0ueVznDfXDmvTPIM7jMxaWQuUUwdHj8xBNbbChLuh3Xf7HygVZHu6jN0dyYXRDctnMAoj9
Jw3K2A7SUh4fb8nBWHQ/K7FZCTrh9vzvvYi3sDLy9nwGfW8mBXq/4VtX80oLyIzikfB7bJHq26vf
6KzoifFGubSOfpnM/CkRu4VbZvrn0ul0ootocWnWAG42GwLf08m2ofiodAOxIngCoN24N1EoRCW3
ncMZUnw7oK40lenLSWrNeryb4aRjoKpHi5WD6tVQyM8e+7Yki9aX4tE/vaallveumpLFYOXPtWdN
FlGoqbxFAi5psgeY84nGFm3VV14CFbwffbHoFhf8GgNQWENVPUmAdilyOVAgkE0Rdsqjc58PXgw0
i32M8Ydfy6t3ne40K3Tz7Nkw8oWyBIGreqrEE7PeRjAPt1FRsDcw90Sh9TYBk3HPJMWEf7iHMd7X
B+iRdLaLaej9Gz9lj6CzV+tHxvvVawk5gwP0fuml4KDrxOgmPiMSQ3Xf6t+xsCMbg5J3V1T6WIc2
smibuV/vvFQD2Il8les0sVP7O6lkwgL7CFXvECpm/1OzRVSDDi7lqIJRX1oGvXePRopXb7/NJMNf
zob4tDPYEj5aYVcXnaIIsFbcO+FN4oGmU7BhoPIb5FV900oFgaKEhspz8iTjvIYxVJYFhR+ZkO2X
EAeSXjLpW8ny7Q0DleIrFW+UItcZHkCStB9vN9UlZnk0hf2uo/qYq1CYKlqd/fAlXt9ocopnsRcz
/oXMssV95zyrDBHGwnVA66BcRSpM9+dsD+PQesuO4B4dK/y6lMbbCj14arWnoz4M+bU9ilL6nq8E
gPSHA8a/ET1+alGvgHbnrdi2l1vwodZ1Ibi5C/pPQxVpwYBN31s2okONevJ2WmcUeCvhq1Sc+K0x
sQqbzfuslCmiPj9C6tkvp6vLWRU5drTZAOv5IfevIohfP7jr6y4GpLpZvnPU2GTSqRDlZr45JF+V
9bsAUEl1PeA5tmKg0t4LvTuNgHu90ZAR62efvllcdCaux3Coz45l3RKZfVEjhCM98s0e7PCmRqJU
sF0Ffcig2W/LANA8rref7Xt+vO9rr9mPL+BzsrysIkKaqbWwbDBRI8jARoEFopuQMhCykbT1ujAC
MrnQteOUg8dR6Kl6NK8yOcWsPN8fENPNxGgRFQx3MtlGKtwLlWv2zijFW6Q7Nj8UO1PYdDqB3KyI
nGTMtmKZTCHyY3NS4YH5gJaofr8SFpBxmwq2ynZK+EpRLBcASNGtcIuyIFcF40R+BR4NTuEndiOZ
MM84nJnfetyPnjoXKweF+B3m5BY9Y827eab2N9tJY/g14ax0SJJx7zh2ZV1ZCqVfqzvmEBvDNfgd
Wv2w8EvU3mo07bAmogv63gI6Puu63FP+KjSUO0pYuBWE78dnF0zNn9+eXbJ2QGtdmU1dxwWwjDYo
MBtTje3vEMS/kOVWOJWDAc/5H/HqDYIPkBUZvSGKP2JVI095dYvgy+8eDEFPQX8wzDuyB2byTAqH
w/ZEq94HOLuM2al5GSjYBuEp3VKSqiAUcJZkjTBy4/zZ0jZ8Jhhl6DPqLXqRVPXEmgUW5AiEZ3ez
QLVoc3Uf3F1DZg96lm7KO2OUgX3IHihoHykCq80kLRXOdOxXQ2uv7zU1IitHHI9yNQfKqeh+gHvW
BWvatXYkQJ5vDMkw/aTxoMV+vrTsS0BMMblH2Ig6yDi5eQdsnTh2HwyZ1GbcYqLgtiw8HJqy4dZC
jrSSOkI1ChnwLg3qUhqwhcZx45Rj9rXZrVzm7H+H6Bb8zbLlDwa+THLb11J/6OtCzw3HcUlSQHq0
8sd78VanScKYoQFQsya4K4auoASsy98HSdNzu4mKI2bLj+L1ieUJGJAI930jpIQ93QR+NugU1oyC
ehl+H55jq7ER4uhZ+yiqBX/Rq9JvqIQHXmvFBqPboqQlfKNCbSjvSA2nSk88BQxjVoLH8YSbegYB
cj4tPKxNTg1yaHuync5C0xUDxr5L0Gj5riKwAOtdbIecvQMAYkZUoX3Vj/7Y3W/Ax7RnvOi08dIM
eHLtBoa+nh5iiJ3AkGTwVkvjSlDhxG7QDMebSgUNHPnScJn02bCv+RJg4dYrbUafPXIo1fRVMZoF
dbwr/v0g56tNenBlKt+Izy/lzQSisdt/gaDzErogRjVzZsH4w+R1uihGx8gzaTifeDfzfwaN/s9U
wnE9KG8gwXXMclSp9qFbtso4/y9QPkPUBjyw7ClxdJQg902VKoUqT1kOpft1cRsWbf4/mdi8WJwf
JqJdBkjftcx0l+tp1Ke8wmamuWAvX7tFB06moYsTvL8kgGa0nW7j9l6uCFMv9HGzfT7g1KvwRfE4
K+w/ABr7bb217i9TMIgU3N+dSjN+BlwLQadAJc05rnL6SyXvGlnC06HdeeugA1DCZRmXZfyjltMA
xBSvLnPsX4+O4AJUj8hTyItcW5ZGoT2ip2e/vbOSxruOsLQjIP4XM18KyIpi0OwbofQCbvmg+ti8
GECpp6exgnuWJisIjL/HCNXfykSY7qQG6rrrmqQoMG3IMGOm+tsd+gtH2Ate5ajd+fIWi07O3SA8
Wr5ZSv9DiayNaYU4scfpAjI7C71ouOmLbQNl8Lr1ywsNiaNpx4E7y5M3gJ59aqEQeDbcgvWpGtPj
VP2tiU9eUTAvVTQWTdBzlEi8d2dLYYt2wjd1ADWfpSBXA1LBVmfbInZ6EdDZlBJd7zs58RKfUn2u
u+VGqosGxLU2goPMFN2tjgsnb7cW2quqoltZBzJ64BZ2x1Kv7Gzi0Jws/LOmNcF/oMg5sXxtiykb
KW4nj4xF953e4ZV2wn1XQaxSSbbUPmv6D9XEpBigSW/MTNTvAe16/BeUnDwxaR1sYRBoBJyIFfrq
Nkqct1DjVkMG/tbMX4F8ikITjf9ur9SM25OGV3Dt3wh6V1q6iGGsYIeXL+/UeUA+M6afg0v6uNAd
GrmZWVITaX8dntw5/s7Q6Ztu0GBInF0baPgtsAPEPSkxQLKlKmYItC9/j6dVuHygJNRwLKFJM6zT
TrdCw1+n/jRl3DIpZRqcI8pGp1S/11tVmWX6i1BHbJ02c4C19LabwqJ3uip7YY6uoJ6S7T9LC9RW
1i7NDPY9M3A9ff/tlMGZPBvOcrldh6QTHRY2aRsdbxYNg+Qgo2WPQ/VopJdQFFSRDGk+Qw2qlcY2
GEn58vA9jTHfgpkv+0YkuaB2s9VMBtnwKIOI0NhFum2Fanvz6soKeDQjhu0oxYmyVIisWel70hER
YNQrO+S4NTtD4w7csrZPcDfAI+oLrVruSqwaN+qEoF6+DAC4ooeEYfGNU7YicVaBlcKMkmBJ/AGV
b7A2V5z7EoMBw7fi6RqvT3Nxo4/Ye6i5i68YENdPKnkjusx3qpJyZSeQK429M7Gx0C5mhNiaWDI9
y90KcacEfOSd3PKrhX9+ktqo6n2mgwo3I0WsZpQ68ozIqIkHETtXcB4EJHUySvqG4DUESW0GB+4u
FtrjSJzuZdi8uVIfrfalLtNXz9s4WBeaYzSbPX6oVLQz2K8R+nT865hG1K0oecC4Wu9uZm55/N5b
TeIYqb7bBwC9Dqoe31uRlr6GwVe0BmDbwNIw4JKW09vqU4jzYwishut2JUwxW7NcFaZdO+RWXwJp
T4ENgYsUXW3HSyNnBXSNqaOb9scKy321bTP5Wi/kJOrLb+SHU9jLYydT0c0UQJ8m2Jlgzb2Q10i9
ENpPDRujCzSQLwQbw+W/moyn8OSr2n63MPKIaoJf4aIP5hILLLuwGD1ndUNi3YbJeyvofH9YSN7k
VydodvZxZmbbX5tbZUQqwQN/pJEaYDX93zFR+7vMnQEHNrb1eXCl32GVjJkZ3Tj7tBX6Ri+Ge0uR
lJtmlDf9gXUiHYNGPelXVRzbllQQFUJjJup3epXEY9G/3+8s2XDim5QQQLw/eV1lQix7ixCPEwCS
PZ+jUGePhdr13dtn0/O9BQMBTkU4E94pA0Ton2R3KykGSZxCxH6rXNP61DomnHPvETdE0ilbCv93
g2C4sEvg3shIhIcnBeHHihFzIHMqiNXEXrr1OdPmf+V4E8U1Ho+BDKd1uFV9IEkRlgtzw1kdZygt
zIrCfmHHF4tegPlt7FD2NainiJd71IkR3/R3KHh3y2I5DUXavVH+HSsA55lgxxiUxRkjqRQOqLGK
7GP0vLmkmbs3C7kS7pvYpzYo8y3OMEWcQIzD8ocxLJsTU+N8B0iuATOQXNTYzw9ZfXYYJnv5QGIj
3LpB0WG0Fgpp5BvBySi3Alrh68KqWz3TLpnxyqgJHXcIKg9ly7TyDPYWJyWL5lh4ZoWBcNYgQ1FD
jqNTAzqFy+aOvT0kNyQdk2iVJeAwf4SN5YmJDGAvHEVWSiyJ2hW8tLnyM9qKwbNkhCAtvSGpaNW1
lWY8ArS/w0QAqcJCDE/BrAjvXd9CwII9/6J/s/i2ltQJod2dsIUCAjzewd07ImZPgDYDLZh480gQ
Q5Eg5P67v27GOAnLwyVVph7rHzeLrieY63hP/38Zxb9v6jZZhNIbrtD+/8m5q+BwOwvxof2Q8/DW
F0VLPSk/tEq4lE/W3ed5fZ8ce2vFOgySmPFtqNBzXFkD3/Tud5g2WIkaVjaI9ykJ6zsCCj4pChxY
iN5OgXhUOSS4G+lIgL1gsZDdkf9Q2YE0kIbxNs4mFxCCy4zNh4+fayxl7+Q51mUXTIiDb9xb+UHR
zF13UNoNiQRafRszOtJEmVaApjVHoKooHNuECgrEDz1nzhGImn1yGeLDyQiK8vk474/u+idDBpY2
oku0NV/0bOnYd4eq2l/hMj6XcPi02vXxSSvMgrMbsURrXAqr/6GpomeUCGGBWmQPp9ezj0yG2t+1
aOnZzRiatVCP/+/a98qTtFGukTy94sHzpAwFEiFnyb7XKD5HA9TwzKq8P+EvhxcvrGFCUHqXssbT
mzpJ6qNbnlamzb7BRLmaw9D8FxJ8U5vz8X8zsmSiz1+6s3gA9rYQXoHM6X6Smv502D5/mVDdZjoa
4/sX/6yD5UJC6wa9BxaeFnx/czyrQ/DGe6BpvAwjWUZDajrjWBYbTw47jb04aFqqCY4xHki/MHOO
u04xjsgCPUCl7MJVLmTsYVh3Sns8FB3X0ysVu5k9Jlu2B2rjgPIziX0gwMQGd+ohiV/4fhXWDmcp
k6WefKJNuUNNyXce4MXr0ZAs+msm6hzhxWS9xZ9SY4NSdTQVgy7uHUbxVwa4wF9SMrjiBEfa05NW
QUlS+P0TdaCsYwQAuIc6LDErQyioNbsVQKZ61khvGZhfzs49HdumTNIaLGdzbkJfuTvjcZXclg4J
LBxOKaDsIBdqI/0pbLB0mhLswEqcM8zWhGv9sH4hZhfZaWG1IJNwuTFLffw8KS8ih9vbisT+Yycv
U1lY589xR5oMQtrHNJJ2l3Vb1c6XwGbVe9pncYnveDa34WaLGJBQLs2CVPef7Y/558ozv53r8D8e
QEHh/B+UV77ej0Rl84SSuxeObJwpFixmnOCemMd0WErTEDAuFgFyhoEpCk1TkUZNtZYZelrhr9aT
5uZu/3hOtRkw0ckgw5FLGUDBoiRaTTFlgwmdZj1bLa+BQG2L8FMDYdqW4f1C4XTgwP7UJ378p4Rm
VUhGRJ8kFrySXY+WvtPKBFAhxlr6H378z3om5dNx3ThV+5xuQ4BFkCaGscwKDskHzjD8R3yw+UbW
ylBdIFv1hV9hYv7K6IiXrGVAh9Y9g9GBpP62cRity7/CqmnovkLok4bMSttRvHmC5CKjagbnSpUy
lljJjST0YSQ6jgXUk9GvK6leJyEhfsf7hsVTT9+60uD6zLjkZtKxhrTy9dsuikehYqY0GajnLonR
aYjlzR6vcTfjZ+USAn94PK8Xv1+XUF/DKB4X+chkDAaLqr4GJaNX8IZomKD0g4rcAnSrUbbw3LXS
F83RYaeshilZO+xjvXN08v6SUb4trdSZiiOTEtmipZYm3HNnSiXmyfic3uMfYGvaGJTqj01k7ptX
bvRw2YCIMzffBqmNlKLXui35s7FUZiOnp3Cq4EWXHb76onMU9v7wagvXBadQBKM/s8kdFx/W6kPw
wDvv55lv1e0pL1jsMXg4u7aiMUbw+AuRtY8d++y5G0WPvq4+7UjW9m86pHePAhMMaJapvcXWnrlC
HMaEJarTkhVahD8d/UYhqiC/Ss45cpA9Gmfl/tCe06RyMYae5oXvSK+f5LhYYGeB2cAGpJVgKBBl
R/RdKpYu5CqhMm+VQPmcxc9+y1/0s2Q+rxlfEPkxMX0ltQWM1jDACsSsYOzgRI93OPcTWXtaB3KO
mRGMryvVMei7DkC7ff7z8F0OaN1khlyD4aHRtEJxokhLB8c+Rt8pIxB3vAfvvs/cAFdyL4N2hCq1
ytu5Hxr12wfxMdle37DkxzX+osGgjDDhctwAbRAb5RZdJubU8v7e8qWkzjL8KhWenzuIngfQ8IOG
55SuUkH8Ia1QVdvPtvxJhXGC97D1xxrqhJXUsBrbv5iKhq3qZFLGjI8dVr2Jwn6yUsic/MMPIuPu
VMi2O99kVgsw7xag+4gGpdkqW5LHrZVtrnuRAFJylHI6zlTJjeD5IgqryxFtGqQphOxnGU/ZRv5h
LMg6iIxs/3Zk0U/ctTy21c6+S0Susi25jo0DwdwO5YX8HbLG0KPR0HW1nm/jyVlQiSgTo/KKa/AA
jbD7I8YGWBFloEoFXVDeONaXjRwYg2SQS2ans+Lu5PYf+VswpVwSUtjWLap2IvQM0OR4WKCCZcGd
Zz53wFqFH2OZZyEh7LfmT+Pf82gZx7xzago2Qb0vET0+MtU+fDg84wkqwIbghw6LOwqh/tYzjHHC
ny66fCH7i0IWbP3Nb4ZkiyNawIfCLzGHTYS9RsoyK4ze7Wez1rSj/jBTv980q36gp3c17HWWh0Y7
VzC2vItA/ELRbGiCxsiBWTVHGuhR0O6SIuiRCMMk13FF+C6qWTMiJ4JR/Ja8ZJdLnN9h4ykjadZF
ySGxL/1PqbCmSnMQw/niV4wMa+Mz101O+pT0NvAbm2HXeuzOLZdzV9ZGlyPubO44URPEw5sMIrFN
g7TJR6tAP2TMrXVVSTe9lMqbxI8ICDqQv28RW1gaCzJHEANzHdA9HmTJ9xQedY81yC2/PiCxhSLk
HWlxa731GeGDekDlvHvh+HYmYwac6cHxeHBcddN8WMwL9aqVxrjTpUx9SiEYj966uWP5qPRceMl8
GC3zJjZMLJqjrj62Ok4jM9IzhQUSHtVcMe3OJvkbNcfyJWBnvvdmUbxrQa7pOKvAaBZNO1MJZ3WD
6l4jl8DCQNbAUY/+gJua4KbCOoncLgn+uabO3Ekt3pjM4W42OO7o4pFGp4jUIU+iXPFs2wIz1M72
3nEaqCutCT4JsEbGsmruxWqRkyfWvGztRrr7WAL0+rwW4g2KfhKpcxl8o9NMq6vDDjcSw0W71WtA
IpIatQ7g0QlSp+2HTqOQAgh0hDVv9lMxiB4BzJ+FVnawQr6MWYha5t2OzirnlLPlAD/Sdkd6CXiP
v4XAHY+QUzStbNxW0FsufQubYBwbyCvUTLjLIAUala9IDe/kEmKbxHpxMj+Q//NmhG7Wf3u+gY5k
zHLHgd+Pwsu9ct1HdnBW8jDynfx0+6QwD2JvgS4gjgqgP4l69Qoo7OioqdICefElLFM4ZokQj2hj
4GyfjXxD7cYFRPS7YXxQoYur2eQ8/q0GckZoZACyKeXhD3fHR824LFLYfcYePzloOetwhwEAtgUH
y253uT3orgHW8CfQJZK8Z2XTd7L7/CIuVpMObOHrS2eAdESGcZuwnOFbnZ7cf+xenPcfFAgA0Th8
9oHxSC20ulIsiUL3DClcNO1gTrJCTbUsGmOJ8DA7iWX0p2o4QdIJa0xnhMyl54trqHFiOITI9d/9
aWPYiyLKARxhcjkNbTGKf4IYtRGuQ1l0Kie1Vnnm2O7cnvU1+UrHe6uilOkTQAyp9vSaPQRP7WqG
NG2dSRiasViD623ga3PSHaIbTHN+t+o4SzXcR/lKj1HuM7GpFpz/txFLVHYrfWofYmZCOLLyAsTn
z81DHukw+hzm5ed3i7l+mNU9sn4Pyjj1nEIERGX43KZ4ctVe3HTstwWYRm+sQyt6QCCsr8iE1AYD
0meT7KCY+mo0jVOXkrcfIEuyCj5V+dF/oQdjcRAtUzXVZNG0WApnbU61D07UXdeZVTB5HcJze8Qm
MJfzX3ru7rbOSLsFAUrH4AGX3wLQE+ev7sVBvpAjg/PLTB8P7Qn/fR70FWY8KHF9CpF1xFbYTD62
U48T8fRdl9mFg50OvmR0PTuy5KnO8p5Ecvu4l6XyJyIQPrWVaGzk7cvwSAM5SsjHP1krEwq/oaE9
mwe6HAZUWL5fCpkziayEpAlrOEi8tg5jUiP3FOo8e+qTx0z2T7kvq6g0N7a2PLfL7NoEVrRSKoFv
LXvKRJiJOsu974AoyFHA8ryAAybotpt0qBxuiocbyJv91DBX1pQwzgOqgeAoO/KXgdr+blWAaLkY
WEn6h9xn6t7aybWIUkbhibz43Y0Gc6TRyPixjkXBZ1a5RX8EfCwfO9LrCq4eK/dV4MzbqQ+j7rYZ
Ro5aSaBQmsGCLspk6F7eVyRM/Neyzn0U1S6vXuk97AGsrVJRTZE9JdqmehzKqNqnh0b63kqQwtRN
aGT2IGoe4VnS23FMyKZodPzSz0/HyzrRzm50lcMjQ0A9HUJEzBmSosXbhvIe/6zlJSstpNaBPeFE
7jCc45c6tPuH2mxew73LLOvw/Ly4Vy2pPe6wdQsCGy2ZbZ+sS/PeduLITVIJ6PsxJpSeTFNa2YtC
pi/HjbOkxLH57nbQNAQaVoZZRyHxngVNUai4EnZorxAKMnJtrQO1RzlCAN0YOtfFilbydgabpSkU
OH5Qf8+l4AMAn369FPkzyjbTl8gbplLI3E3w/wGQ8ODS2DlWrp3EmdO+RHcpTPiMmMQ50K2UoYSY
J+9hrl2w3wNLDzlnCs+lu4hfqKg+pfVHsLN5Lzy+4qxSlCxiSu66B2PFwHmh5W1FudSLvou+rZvE
ofPwNZi78Mgg5u4HD7dCXKH94K+dzqMfvkvLdC0fTkpZXicuZvOiyAHYbysRtsZLgyu3B4FBmguR
vW4dnd77p2UkH4uIfmVC8b7oYV9ipizAzWngBT78q8730qcIkWYmos2hcbOT1Q/zX6Jguf16v4VC
f8SSXjwchzEV3BCucSTqny6srQvMwl148qkmpOcNopx6CtyhcCgsimMdSFFwkjLNlUFcMfX+qf8v
QVWfxOhRryxB4UH41eud2mmIZyuq88d912Hb6y7G9QroEmTEvzApBOisEu/4icTq9W4DUNait4fG
ZmDn0UkWMyEmKFtaTkvXLJxbQKH4QimkRUgfOYwvH9+APIn1n1HQNkIO0XWrf48BBCgEbDeue6RJ
X6chLSyReqUnrZV2lHzVtU4dMv/EGRO0EGGHgCXuKpJSyVHUlX3UVx+KtN6xYnvCuruRv7xR9Jyq
G8TfRfQMnFMPVSjQtEW34A+xontMJwdiwmCb129jacLRNMeR+hbXSJuyRPuYkX1YSZvPwsqMA1KO
HMaq5Oq6t2Gnu8aYbGhlstAE9HrZZ2F2uML+Yxk4vIazrTagUMpBssXtP8E2GXsgmSGovfzE/acO
/SZ+/Pg+sMxNuLyfIJz82dc/LJhSpTymW3tp6P9mtyuwtNgIc1swDqmt4DHD1nC4lgs9uQpOZ83M
I89VsUpGqia/GILIqXHK9mwdaFn7N6hfPV+MzlqVmVMtncx3Rj+UyEO2/uVAh55xh1Qo1RVxEMlj
5o6Nh97wamDq52s0KoMF5rjOBQecl2guE099nxDN9AriSAIqGNPIoYt62vg+VxLXCUzsSa4AXUeX
FmxdHi2zVQmaTQtXPuYHjfg2V/aMvAPJIM/a482+03dh+NGMpZZ0NaCAMz7m1E+BLTE7+OPyhfT2
R9epo5EI2P3nYA+Y2ixBjgB+x6ibcBcfPvJFqO83iwXS1inTOwWrGyMfW+R4Epj0kA0YuyT1TC42
dP+E6UR/JzWfd57Acv/Zeg3aeyl5/9caUHUlJ/dXfJC0Opxg3YVni5Ng9ptuPWg2s9GNdGCZKJyQ
jstjbZUiV39me1hFQGrZVxf0sMMrBMocPkLzZcaxzZVrT4/pl7WVWYXnOp/aSUajZQ5JKCOK8D7o
DwbNbVAoT8ZScUHZ0vQGHpn2r1GZM3I8z5iMIybuTXqsOXthcm0CJAWPMTGKk9mUh4gQ6/mIx2g5
BMh3xm3uQiBHIq9w32ktZfpBgltn3fqKLV6aFLXHTB5Dk0gp2dw/0B7BXwz1ZV77dfnsQJV0ykFj
T9VJvHQz60ee7mZdf+mn14ew6SmjR+blas/YJE04dFfiuYaZLd0QqitxD7u/R+2dDEZfBIlz81nt
JVevsZVK+46Z8RjPtRb0WBklS5mXIYIDliktfP+cdeeoqEHmeIcjr0bCh/lRCAyNEtpaoo1hNEAj
PW2RzZdnOl+kxJv78CTQuKkxd5dYLKT8MH6BUF3sqh1mnBg+5puoZnMClYZ1LC/7lXTjaeqazeP+
X3Zj8bwBbTVu5+BEptfJwtFFRmK+YX2VgxDXVry16gTd4Ac09lQ0Lz7H6YXncdh0f9E8C9NgJjpo
OoMxZ8jGdaSTZ0ZNP/CZL9EBDp5qc9rSDvp+9rFJWMtq91JKI9MRS/giHRWRSzlNG3PG4ZsG0zqe
+NlpP92UnyMoThWnjuOcQ2qnPJiF4p8EgflU8kQx03tD+NP2OT/FtLrSXqgMkbiAhYfcrnjC6qQS
gFWjWw/FDUJpYoJr3rg1FE/AC5VXzYOuxI+1t/GQpiu7cI62q/YUxHqO688gPKQGaLtdd5E8Q6BG
u5TpA0zsF9DgIZsrkMRbgUEaVJapTTt5D3j0OISRuSL8+43//FvFDE8FQCkuXCGTSUubo2eu9v47
eCcbjD1sOtV2KuwC67W2NPu/qvPHr2koMMeOhizvgEAapvDroAvaZA2AQP1kT5z4E+J1Jp/+j5Nh
uVdMj62piodKos8ghhL94cGLYvtEoQ3BERSl5Y7stA6SvO6OshN+vyaGPTIOC8XrvMf0AmN2kZN7
OM+DJFV+7uTdWOXV27WBumsfVtS0x6Vt0Rg7syf/p6FRqSJ8i1e8MyapmRKXBw3Qm3Np5I4Hp/rZ
oLf26KZoHzkXaZN1Buh8ra/ae+Hxg+bAY6tEhLOIkC6IXMRSq6HcB78U+FiaLEhmE56Qyvlcagd2
o8GU0VUmKXKApcx+iWCBebMZBA9M5aJ96yF9WLGdq+6Kn3mNMm0ZoCGAkn+8rB6nKtJlG5yrkzan
xnlWUO5VrahFP83ToGenv7e/MJ8CLbvz6dhCy2yQxht3oCAhujs+3jbqBY3kjO/Subs9yZF6FKIw
nSnNqJpTGGVjs1I+vUm5+7Hg7f//3epEYYJ7ptyU6BQ0cxoCR0XuolsyZjQb+dF5I3gMmmdrZ4jG
/xP6BtoxjDRmfCSXW7FYTt+R4b/aPngYssX7gHVbrGHQ6ZT4+I71R7rMUN+45hlMYoon9OU8Rc1E
frZzYFa61D35C8aGsIOIoYKGzq6D4c280nhu6TqkqweGSXKfvXaJ0mxG2uQ2X6e/zGKwk6dqshIf
MwUtV7JOAST+l8Arm8UIV+P//MHuNJ1AdNmrqbNboDgyopNdFIjyLz9md+RE4Jq4TAz8yUhq8CJc
HAPUAPGkmpMyEpkAGgpZPf+GO8gEixeyOAJTyzeoGyMucyHGXSKNZ2hzdLl3UlHAgGTUh9uf0S4B
gCOYQHSxsKmgasuXtPGahbQUf4Iq0+Iulp0gfWPr9spTi8Z1QYjmZMDLqr+1HySqrBDyGu0xrPcK
QbZ4MhOp8/3ZH777N1eLxR9pIvbOZMGNSqUbGVUq5DFOWXR+mcxGQ632oKKDIEy0a7TObWZa3GSi
rau9MWH3LCIRnfr33+wKebfupaC0K6xpjAKFovk52sdspKnJz/2+a3vCT4ubx4L7Guu6m5lTDMD+
g0iKyxWsCUwqMYgQGrXYpOhW+s7ndyluBonQ2zVvn5mhcwtVpiE+VbEAGIb1X8wld9yDxnv3OLy+
BKVPymNmFWWXe1dl73ZrgP1MPUk5qF4f8At6szZ9J0V61rIwY9KTsq3k7o6Ds3dq/uv0ImHy15XQ
5b1j3xgXvH/0wTzUmaHB6vtPY4SncwkKMI0dMV3e//G2WEiRFtDjQrScIcV1JI8mSFB8Bzwhn3Xz
nTTrMOjZAlzvAnak/jEmXwJkLNLSMZ4vLWUNJ15WnRb3H+aRASPB2fvmWSiy01nlsX44Qhi3Ik6p
apQTkt+ZwUuvcETsKSKiLMm0/3AyPJLv76lYy9ipjjLUj1H4A3zEq7zk9Hu5dTWSt3yuN+M80cCG
Gk36Qmvm1y4NGm5OxZTFM14rwenBFe+QGiN7z94+NYI/MSnGDoaunbJc8PPASnKln6NNgkiz2Qdn
cWkpF9KxuJh3mR6ZBwbTsr3r3Cb7BLY49eKf3tR1LLOZt54m/HbxKsdot5tQIJ+teUYkj7+G6hu4
EgytvP14m8Lf92DLL0U+VWFflUqJL3Xkq2/cFdzrsQbYlpN4UjFS7YSJzlwP5BSum6ZMbErcEmHv
w94jZWi7vUb7jshj2nMDn2qxjnvKmilYF6OUiHiKoxg/HW8VvwYdvzcGjwWZGRt26K4gd42QfcXy
3VfqZQfNa97ohEvgU/4RP4Ue9VspoVBc7ltU/fgRtkVnRrzWLNBPofb6eXflqUvqnKCV/6wBt3Lc
piuOZwp+2SrNvOi5L+2lDLD02T32iP7wFqSj4OATsLUrbgm5eP5UJebEMlOaYZ7uZCDHvy330h8O
pzhMPTdX3X8tfKw5M/9aKH+em/x3cQfmEALXBXrCgp7L5JItyasMxJAfCVxDJ/uhrxQRWoBN3BxT
OeXxmSgEJdkeAW2bONrK+t3rdkc5o9IOW8E8SIayJH/QLzHOaiNv5dynmNRJtgxFifI4zzyX53lr
pzylsBydHzLgzEExt3Kyr0nvM/vRGjwxPbtxwuelfbkbrcxUMnWdfg3qFiK4mFUhu27HkzCD981s
XqBBZPewoN8MtKi6ioHvh99pm/hLgfhQKz22mMKCio2VTG7gJnxyysRoixtO/557x2DBzM37hT4F
bhDCvq3ZnnRssvre0WLjPqYtN/YDqr8Haw6H8oGnUBa9q6r3qR/t/W7QQled0Iy7/Fijhh7daGJd
/YCSzbM3dPviRNMDqMY5Wt7OtqOwV5Y96ZJhKKSVjjF1dpF7zsbcUuq0IEVzcIBfDnVEwVsa0TqV
4V8nhE3UkE5PVFxDbGG9J784QXFP0T4VjPkKPPamh1fdIH1ik0g+A41fxn0FCoDQtsDovHr+Bzsy
mLEEstfnUjIEzRhi8H0Snm27JAFpDCjQhdQPEFuGOT1Bs/foNtDgylMbYhKHMqtPPEDmy+pxZoEI
Sj06bgM0V7A64QmINfv4rb0Xs5MpP9cm5dd3h76MXnktoa+Ngr53p4GCqyh2lA/kdQf7ka8yZqsg
jIk5nbp5XJi4l8zavv8pq3YJIeBvKGPwwiIxjWR8ykwQMIziPvW7Dsy+/KJEaHt1t4ObOOn5ZNCk
ZKjhbaZq6ZixrujpoOC/fKZFSnh6WW6a3h6R2ErVSNzgYCMJHAY2GJOg3PgobvP1IHGAl0l1wIEz
Pxal+o1PN6PNTxeccA5VUDSiyNuuqXz58WnZgFe1nhvRQYX3zNZixNjcD/QfaAoBWuTPllxU7Q4n
hocMVFisLWMUMUNJF/+a9wPHwNb7g953IBWppfPibVt8TG6AEzGF828qoDLx5LL8vd7zFdB/Aty1
t5cXfWMOw7XfFMJFGPHmuRLGbQpGx+ZLbqrYp0nL9iKjwF/9f8BbzFErbhBuagyUTh1yOoJanLL5
scJi3q/8BQIAHRj7gY1iHPVuaCuPs9rbxVvCcovAzG2RCrzmgAaZJ74z7Rs5Oz8rQ5kl1GOkFEm5
gIOsivnJ5vdTbl3sPxejJDzT7+zUyKc3Cp0arODQppd7gF7qyKNJ00MeIlyoXAnw3Li6REhZ1fkk
Lr4BFGxJQqDYTuaihgjvB16dr9M/YEgDvqH6yrTFW99UTLo0n5DhLSNKwg3qymwvdhEgifOrnlUN
8VACipBD5pMXwdbiiSjghxgnVD0EKNIR7oxbovoCwJ8lwsbpExXfVYJK1YmxNn+Zf63whoP36/yH
Z+dRhICQqyQwbKgE7t2QWsz4g4weDA+tiVTL4PeZgPQgts8P3Qi0/ncVvmw75jdshCuVwexj1uHr
vDi+u93IBKdYMxKrA3pdLl6iK6ZRoS0yUFd3E98UjFhyi9zybva+4WyGfgtQa63qMzQL1DIrfqLz
NV76O5TwNIAs9Nb1Bd5JWl6xDQyAkLbixv4Tp9Db+/RTyCR72cPsRNpGy2rNDJn6E8x4KJlZWPmu
QbhIvv1JU7IqOsRxt7+yU8PB2UPV9qxZrVkEN1LavTw3QID25V3BqeRpDhR9a9pW56QIeVJs4BhK
nUYSJUUwXFmGVA82RMM61Q8OWX0yXJoZ6LZYEKNdOqQO2HXiqhiw4G8qo53KBeW0VgqD91M9ui4Z
g60IWaG4noW84SCFbjzCvDV8j0QHVpQiKq/iY3GBWntt9nfznieeG/sPo/r90oxed1tsqA24GJWi
Ua6aBlH1wJ/rvab5NPmOLHuzHCtfMdp/8aMKED0o28siK+6rnb0bmZlzLzcHsSA76kldF7lX+aq7
Gub0wlqlG7n/Swvw+psV1H1SMinyZEfa2IW61AezRq46AilzM8IHy6jLrrA8TPgl6PtQ/8+xFgth
Fr9cE89CleJa11P5O83MNiWstPQGDp8BlhmbGnXUAIPwARNfpG/1HUmZf+33o7XwEADSNpzpOBEb
tofRYJBG86XWiQk/c/EhhCc7nC+TTldc32KvnUn5tZ+7Ec1Piy8EhQtTUiocke2u1DpUy8gbcfL5
e/HeC3iHv1EazVXa4PXiGp+Ty2zveCiV4onNobjU6Ar7Q1r1Ria2+ry3wk3nn1cyyG2WpHKXtBH4
UNZMwxt8lIygBGWjIn6wh49p6k991oxFJTF2o9RaqqTYh9CC8Qe8Xy1oMCjEo6TtEWpljO2j4DQl
FsShB3EzPFoj35y68AuBq8mTvpEpxi+r0Mt/YOd1PL2AWxIyQjjKK+060MZN29P7QgLsA3l4kkBC
RtKizQTSUoLY+FX1zfj2H5a6R2d50GmN+ON3xqqHa4kBkQ7gZy8smIJcLRJryDvk0N00s8NsbZp1
vrK85k/bPfbdcsh/9YTflvO4gJS1tPkDcgbUJqaWMGUgcPbC0eJKBQFP1N5ii9tO2+wovmjVIsiy
IgrJeqlyh+WAyIid7qUFzNpqDo9/ryx1O8Zj76OcmRzrvO01qqgsi4GXTaGvYUBxPo8ohetya0aQ
BNOCET1TdEpTKQ9JIEZKT50JIGuWvDx8Za97KpJq5PU6bz7Pio057NsnWPXw/UcC5hCrkOGGs+DE
BPWtYvv4fQAkemYJ9TyQgOgA17063JmOkzD0WxsBzvxI87aYpCULo+57Kmk+hQa3zSMpAiegMWYp
Il3PSbZ3uKLopP3LwhsO02X93TU3kik9V3zpgynyDeFKpOav4itBmUiF1yuHfv8Y9A8/Y5f9NBV0
f/54trVF6CAFG8M6lbec7hJ+JvKBc36WoNWgG+ibu2NAF70t80RXacM8ZgjomIaK7qTrnGaxz/uS
iURC4QCi4W5H8Gzrcgv2VXhJa+/1hieS9tJutUAW2M6u8D8MUihA/unPtduS48fSrhwPd8O57BDp
1nMP/TKnuTS5vpas6wW65MOGSczcgC2pd1x7pZRJGa0z2SYKHK1Ab3g35ucRAHsWZKYiymlvzG4T
bYTdXzCF5fNFNHQn7CNtGoCqzOhRIDKMQMX9tuRoiNT7d9cZR+d61eNAhwiE92wTTdX6ShsrZmk7
yulxgJVPOqVJV4uk07CNU6Q8Oa5A8wPezQ6cvfrelhtl9RXav6IPVYHEa4QLJ+oWenjgG9+XwDZg
JKMGoAsMcboZdyWc6IItH1v9PwnvR+sfBhxG91dmtGkeRwYdbdHBHht4WdUHYjxLyzOYLQoGwKGJ
w9VbUnz5D2IuQtH9rSCOw6fNvFBc/KUkK2u6vy1SFfW9Pya5GrP26vBBc6zQ5ssrckcOhcdEekGo
YfQ1lhHdIWHTMcwckWwmMeP/ztCt1TPnWNcEAdugct1n/O03XVfD20Fp+BExDrWiVyDZnpraOECB
Gq19fSo9Cmf6vEmOPeWsuunUP6B0vB5zdvJdqWK5dnx+yxJxeyqOVLEWbF13TS2AE1M3vi04EfV1
uHjVZLOb1acIWZPyHOnySQujff9cl3vaIQxIyac991ipUztrga6CGBAPuEeIp40NQ5CIEihvhj/8
PEeuI5MVpv39PWuCILEnh8JKqfTBJQaPdH29DcLwSPl/AuPR4aLpM/Asnq+wIfeYZulqJ6UTqVwn
nmmLMS9M/BWzR2hxMd1xJCK/yvis3Y1gJBfb8aZeeCTZpGPzIaGnbib2/E9yoeujvibFjAHByojv
vHW9Jggmo+g7NCeAN1W7MJQxT78ExpK0tLJWWLum0FjNv16RDK4m7qnJdfKYMwEUDSv/x7PCym+2
sdMYWjDTeLle9sm/4s3SwnCoDq2s8JafcQIZjy4ITCbwLiiy7B6owxfkTfhKvvrVHmkRkPxnUjl5
WZ7vl6cAYnwQgSdzqy3Vi+xEiNYr6Pc/bJ4jbegIzUWqRYKcHwE+5FnOMKocdDiivdg9AsrJBMDx
EqFsdlXseQtNtlGBlG7eUTlgyTc6nm/TixuHiDBiwj6lFbUI3qw5B2JPr90RlAe1o67vtml689ZB
cWVXInHL37wjg1Oq+U/wJ0wRmP6ElLXHiPUgMAx9lkbg/IcxjkoGaWNU411Kkx9Z/V+z9RKi8G7y
WyzGcT/mtT2/+DXJ8gu1ksbIP6x52ucXUPITrRh8r1XvZb8PY7z+IAaJ+8aLrfgsOqhUvAvTHzuD
aVW4HbwPApqk1HWd/cJrQYVYuCssOSvByT9rCOp4a1pP3TGUEU/fjPT7d3VKpvpmrY+pw04NagR9
Zdg5wqE2P8kRFMeDOPZJoB5dIw0MgEdONDZhlgCS2QmY80T09OT8U60lAPXiSoCe8gBBy+2g/rBb
z1nPr4h5JxubzYtimCRqtM7BzoXBVazM2TI96kS/f1nNZrLZmY4xz0W0BfG4hfdjfO6CQD2jtPhC
fVu0Ay70Nd8hDjVEnfYGsOXYTjJA0NjecT/wuNAoKkWJNvkICESDrsudet5bgDs1p3jCMJeg1eH3
GM1W24xhFSuh1ClpoO/cmpK3CX0LS8r6iHhUnC3Fd/ITLlWBn+m+wfhG2IVzYrEMQCHiDGNh1dU+
4WULp0POuCfR7HUKtjgZL6i7xYKegUGn1wjAc38EaGjqdjcULxUbOhAB9vSYPUW7v5Kqk2IzcsjS
9eotiSoEBgRTa2izgxmF5wbWodqhABxuka6JhnX/PQ60jiimvmCxSlXe1Y0n79KXCnAHQ06umfIL
rLqrXPFBQkGjdUexxapZYcpxNLcuZspc0/DKqLTL98v91LxOlOOn7eixb3R6FMQokY2DrmM1MJP0
meImFdZ0vIeYe392hZK38lrdzDUmSvI9nnatfKHc7iDEzrCgmOMdXDgOVRMhufyFz7Ub19TSMYlZ
Kqu0B3HaPVbyYOm1yF86Mg3E51xoojDHMKJaktuV+7dd10oS5JpSk15J165WMA/OB7nLgpF4F1k2
3BzRmr28iV96jblM/qCo3RJO6lUi1jtQ/S7VsV0i4OIHO0YTDmLnpCqHZdfHx/PrdSRRWqYRRxMg
/GjWw9Nu10SNdgaB+XcXW0dUwf+KDETvFHqAYN3HpoYBjJ6E5110pvBix9CA5x9XG6/8SDz5Q7Pt
Az/0akrDnK8otusGELT/FltPFQNZSoe0s2B28usxSIfRhCZ930j02e6ysPJOly53JjBe1nVJzkrU
H9lQXW0Umh0txZ5j8+g8Rq22G7X5Tu4MfCnkOwpyBglGJ1mNFjfkzyQsUt+YleLQjG0GjjUkquu+
AMPP9KLaoUvoDM5WhcyVIctQnGeU6wUTUP4amBs7d8dFC/y/X2Io3H6p/UUjxA674wLvLJDSM4bL
LvAMoi1lJjxmi5aCOq505epGuy+E6uZK0MtUhSc02RXuYV/Eb7sLYQt9lyK0sEeQtGn678AvNpF9
1Pg9RQhACGFLxAWCUwma7CXNAKqafK69iH/O82uFA2HVGva9Yw+gxCtfTHO0JahbOxhZEF+gyb9u
nZHg6CrEfw3Eid1kiL/LUO59eDraU93qw5TmsKDkRUxnW8yKhjnvEoentXWPWwgxz68W9wcePiYF
TjEsBYECWPQSvgYHFqczzzb2FmbqwAwkMJVA9JY32afx/CS9SxK3FdhKRP3EWzSII6w8+NnrlVV+
5/0D2IhsIsJ2CwGWEfECvugDqdVkFrM0e29yPeI+n9EhfZECxof1wmba02zAloZzAo269XPL3uuN
z+IQWH8V6v48n54khx5YiBM9AnnoWPU8MxUrsmSityp7vQquA/Quiak2NK3A1YJFbIM+W1Xy7A8A
omKzl+txqSF79TpyrM4zyKTJzvyVbzuRF0zzn+JUHiCUX/unWOeOVBS+vmYOrzLo7mX0tdiZfsXh
q0DuMVnVYbRzXIC6BWcvTpfD4u7TVkD0laZVESCnNoZexNpglCP/QEu9HcY3fij3z59Sa+iJ2ZYA
aY1zmv74V6nt2ey5snr0eRcAE7NPEXAPayUZlvuMdflR4ql7rBiHUUtCmsLSRnPi19T9892n6VsC
5XQJFBpmWKujreT+dTXD92hf1C1CA4NXAU16xf95OkOSPBz0+ovvz+rTYay7pSME9DyBDjN5U0J2
ZBfwgXRnlM+iMDyBY3/fVEE72hX+qw5aFyXhpSWbaKWMOYqySa9dC5IdyKGhXXPNhtlk91NXtbuK
F76JU+wn8SCsqnWxNIVhuwKxPCrlWUomgwCMpNn6jnG9e2MirT5zTvtcXc4497+zJh+rclszxZKp
9R2untMcSDO2DufH7nToJNGdihyNGG0SgcLxJChUAhgYwuL8zGOtY+vdBMZpc/ZuxuJ6rIo5vDlw
lL5J1GgnMuZXt5pFP61CA+OzUXQjxBqd3bwgzOR9LH2gdY3PWUTsX/Ypx9WzSMkKM6+KozBMB/vh
SPZhIKiYZg4uW7n/wRBvFiJ/bbHol1Owut8+dR0JnnCKNJILFzErrPZLNNZdtGBS4SKVqO/IDgb7
sIBWK9ttwtTynKnrIibrd2xm4x9alNycXoMBP83H/jX0nt9+5CmkLKcG1AFfHi5j+0SVw484gOK0
/JSvO2/wc4LGtAGBJB9J8TJ/6LRslYAiVEvJ5eA/3zzL0a74DoFTuif7MA+95LDHFrrPJYgJ4Zmm
2ogjY4cqR8WkX9l2B76YfWjN+zbJqZksbqTUCcanvx3amUz01zq+PpG0uEg3+TAR2zXQmOEoxJrp
H2w0V4CSTLOHX68X+TZXng0iLCBJ0prXsoxrx28P3uTs37Xo0B9EwpNgH2a0Bq5JXmGi5QZ3cMNd
Wll5a0GqlgmmQsC5A18QGNUiPDYBj98FLMMxd1OnfX8BZ05GMu/Nu2CdZOm9C7JouOdxhOVvkGFb
n5qJ3eeU9mJvmdclXtrh7TnAHEO+myJecMBAwJja3gbInfmKITWLtxMSk+jsbGyZcU2t1+RPrpq3
Tjrc79YyU9rzNd7PEJKOgBA30r0ptEy3A3x5q2jEeItofyrTl3J8D9tDtLHbrW9jxQcSb8CH3yAN
8j1aN1lV9T3ooWhgHCzsWv0+36RP8oGuZSKlcEguWEoLTZMSRCvwsPDCCV5BRgCcan052Wu5OK7y
VIzie7x4nNziah4dS7TDwLlqdHN2qQj/jtNdqfRX5r2TmEmt3cknda/3ifVAVXKLCy9DTh5a3O3S
6YPYsNmo2hpHuH287ieU6tGz26azSW+3e3m2hQg48XrTd5xmasv69YYQlVwLv8oCdfu+fBXtO1HM
QQv1aZiy+pbMY24+3Ch20O51grVRM9QhKNW4uF4kPO/VSR34Wn2zXIn082Qc92pn3WkW45xsX86C
up4b/SfjzwvBLX169k16yqY2No3urD5IuNAK9hQ4K9XzPbxQBHSzW2Pjf3lNtNtp044KbCiA6j2x
daF31uflBMCnF8pDWakIh8fWZH2KvwsmVfxgOE9OxT0WxNmOJK5diPHvfiqIiOcuz8axNRsDaST3
qYOcQQ8SVFe+oTmFRJV7Jc6nALy/F4D44aiIOpcDog/j1A5IbJjatI8LVwTubFDG9pTMDmFMETKp
jbjySIvJs3NOb0jniKKxxUN+hSW2dyZJEFyTCKXUM8oI78s8fGVJjnWklMZ6c1iGMh8Y4AekCMvR
/44Y79nctPL4sJ3sfXlic8lohoVBcic6xQKYApKe4PfW0D03HsjBc699M53Gfr1QV/CHulGrhpv4
oIdYUL0lddH1ZQPGOJ8QoRxQ5K/PI9lggmdBv6GtCPgsTE1Fi/077P87D8L+cJi/oVLk4+iA5hpL
1lXxLXt/ktWOJP3ULiBupsjfdglps58bFXVyUIvN9l1UbSLG5HBtgc8K1X+kUrY++MyI9XOLTqnh
h//xqWT5RsO3L4evkxt+nOVQ8FVJzjKVQF55dlOGdaXwEdUY1U7WypCk8e5ulNp/7XEd0JAxQVXn
TwInd9IMqCz2FWBUMyBUwyFRZd8Up3J30b7OCc9ipqXoL3/GuYHVcbYDAG9g7K5YF5Uw6r0HQbm5
LgdaL0Jay8yYulBXE4XGLF4g5I4nIq5MzCb0jIXM4XNjZZnvVAKnYJ+sJbN7rlQ+LrL9i62AZLqN
fc7kIWdsJ87Rl3+wKMkxUUj0+8Y45zfY/5gH7w3G7T+z1mCfRjnom2zl3mTBw1UedST0yP2WcvFH
E0hzFaKfsnzXIz4HHwX4+ljrI/AiQnH9Wh+g8CKrcd7fam4VMwCnD8d3rezpwV3JQOjIyJ4MF2+P
BFeqm5RIRGnB3WCqaDV7gJg5BQfSxvni8qSUmdBwWBSmzr3trKsFNmr/eDyVDe2d+U+X9jFzuYV3
CvoSg9BfNs414TCvpy+Sg+VYDdcrqMtd+NxMv8zmPBqvoLOwCLNnozL7tPNPTzDKgAb75IfspZWN
WcLN3wqAu+cGDUm61FgZynaQ3uVIdoDqgKO4swttA3Ae/gryxnILyfrW4lHFN7+XZeHGPJUD2kr9
I6QemQDqpB2Aj9WV8t8Kmj+XmYOTGTlimhnocHgPlZlyEQzYc1ff5cae6VH+p4QtS5wxItaxdP20
aQ2rkzpNest8qvvfjoRCmI2PI4Z3d+obSWR5rtiI6R9/e8cSbEqsr/Pwm+PqZDRalxv8Ta/Cy7/Y
Ms8NsQuI9CF4jxm0etl1zT6CZzo+mY0cD0UzFqtlYPywox3yZ6JBx5MYCxWmJVUPydDkN44i7rEw
ttMjeSQCt4j51UIbdhJOi0XnpZ6VusFNJ/e29RTbdEs/zWpISjb8CxO2fAEP2tOF279K9KiOAg31
G0+DVxxgP2vG4Lo83JGSo/iwklHHTu4AuihxubSWrjGo14M+qaGd7VXTc23GITdxEk8uiLnfTgH8
t0/Bj+Z1NahuhLR72ihnYXZJ+g8p5gZaWVMhEIpon6Dsq1LM3qGirjLrvPheLNXCDZ/tJ2v32Cau
nUqQ3jJtQABfMRnyJOfitQelV27kqRjLU4kv0H0Trva69jwGSXu4q6EBvqL/ff3Pkln+QcGaq/sG
sia4QulaYFzl8ptPuyLyFrdYMJ3DkU0/ZIg9kdoQ3HJbS+wFvdTbzj1KRqnGX9oR1UQNDHPsukgl
kCk1p457nGtUkBcZh3Egb3sXRzvYImqrqZo7Ch82p0Htcj2MMtz2o4EMFwgBxTngzx9XqrjazL9p
8zy3VpYs4kMMNWZsowppS1ysPD9omC93SArMEOUa7xy7pZW91H1DR7MJX0veaiMdwFjd2Lct3pGC
XumzTbsSpFdKcRcrCTgpszi83mFhFCKGokOEnb1Bgp1ZfQCn0FQwwA7R3EMpWu94XEOj/JWOUROm
6JP+VRocXMbXQDIyJUNeB0YlnyORclcIYaLVMpXCpOKAzY4dB+M6s8E3bycoh6wPFE7yXvCjv6P6
vY2vdgjBxueZYny1xenGSoEnpj2bBWadAAl1jBFC60ULZp0YZh4Eyjglq06rWE7yfSigI2Zaoqcg
3v2Q8x1hnjppHqviuAYXcT+fAcTdEIcO6UAdgQ9xQG34uN4G57kGcjLcr68YD7PYdu04zrgXhxCg
vIC64DpJ2aOOKFXk/zi5T/fILcZkAKHGfu9o3BmR7Igv/8jhbPA6uNTh6LhVUBXp7DQDZekdbVws
aZv7MHR0xXZJjV5Bew8itWCBUz5ZMCrzYAAFWgkmbnWQ5wdRjiFGbWL5CRsFC9zk7zHvp0RAlPsq
gIkMs02kthTFTgUNSHEWxtlnhzY3/Q/xyTvFASupMoUUh6I+1TaiC3P60I2vDih89MpeKB+A6gTE
FB5m3fzVfutnLf0ORcxzmINzg6r0U8wPY1Rspy8zLX2cmSjDz7nsBT6TBcnNKvXH0WGBtun+9j6V
lyBR2SV5oY8HIV+lCvqb31jz7gPwRBo2aLQrWtB4HQJuLCKEy8qENqlGnkH+eP5zK1ObqCB52SdD
saWeMfssS6VI3Fg21wxPfh97+W2c9mFNsHL6UezhiFtDwBvRnzIGnSHB/qw4VZrBZeXTsw3bPClr
H3JD9ggN/ZvU2eWFSK4ePj3Mcw23L3Itq4HWhjmIk5GJmN+Yl5Yd0kDZwq20OLEH1ZyiOkJ38EdF
qcrkVvf3osnu4yGRdXLKsA2j7vChzjZ1nmBcYeouLVT1z9/P7ZsaF8rSFtVCabNv4uZzJV8UVETk
7z9WBudy0roMXZdqKtBmM62tSuBOtNd/3NHggkLtszZP1MU6rtiFZ4n1zqWveQ/neKQcEwHZhlg2
xtYQ0lehPr2XWUrtl/FFGST4u7N8a7x0uh3Wxk3yckQaaqIoSqwH/ZGM6k1YYFQkNtC7jxjNWhPS
zjRDt+kDzym/UllFEKFB0lfTmQD7T3TW1hDpL5LSixsnHe6joCryiw7Ga1jj/Z60BD2RLm+SuWdE
FQY1NkW6EqHAa89nCg7b2quDqLst1AYRs4Zfl3w8MxGM5wYVyXbpQb8FZeX7JAP8VvYvm2/NWXIL
H4e5W9GD2xA17Kc51MwTJMeWaZNnMq0rKNRALcQGveFJvP0fh3XK/fMV+CHg6+YWSwoJfxZL6LCB
/ElkowqbgXsCIkfLnouI0rahynyQMclaPDgzMvbpYa5nMnqU9k9EqBLhbKBz+Og58SzJ7XWLMl4k
8to4z3wKgDFcW0ifFHTiiPdDhsuYRAdjVLNL4DpteAIFtRlHYYm9JKocany+8DttHBwSqET/Z7IF
UbGr0C7d8p6Y5BZjp5/YwO5rRN91re3S9/be8pu2dsINH4nYETMhidY7qm20oTw/weIX79Gn7Gt+
zgZKe4317xbYQhBgJDEqRU/aNWEXwePInfcSAKn3/aAG6q7R3F+pjR2LO/lHx6cJe05ORCq7HD+Z
vIDw65Y4fhb+e/m/NmRsmRVeEabgH9emtHwWzWqELbof/Wlj7zONUyIjFDV94KZlAJN/eL9n2M28
tl3Msb+P97Fclsj8ELWC9QNmW4LxHGIU4Z3Mppr3Y9LDIEIJGAmUFhNIRd1swyv0JvHBEMwuPvIq
9DHLzPVbG+P5SiXAa/QVqKbZhXt8OuzhJdxqTsr6xQQVlzzPVtyHiSdLUOp5vNtzLEdEijMxelJJ
v348dbfJctZVeQoi0ycviT+Gh7/+yhtgXYoCady7erlvZpekXp1arwG119lzu7RMkTwyegIGoMTd
Idy5pUREEntpsgjv/y4fWJ7KtMW0zD8fExnwGSQqMufK/45/qkbUetO90/d4ywWvRLPFHX6Usd35
c/TjlRhBQ1NKpCdZVNyWZxsgiXpR4qyE5ca8m7Mb8FjDTofYLQh9dklNQrlIFDMUaAXGt93O9BU6
4y3sGvRGniw+P/P9qsXw0STQSzWsaTCWehteXi8FQ3mdEWdkFPKi3Qg430MeQ0KOr2d+WLQTIct8
BDaBNHt2tYiaVWjvk+ipkO+SVo8MeYuWcJqVei840qMJqnqZdTuzcX8UaMmATXHQKL3rXHRyGie2
XfieKKS06Q9Xd24IJhcY06cPXJif3WrkFnm9T1wv5wZH5OwZBV/6Idmks3KX1WNv7NDib5ZO+vao
ueM5/HimulvBVRZ0SUVLumzOSfPqh4RLsh2DHObAyzPhw0jwqK+FtznZhaK3OqfktyEO7TN8nhtD
TqYznRfccuN+PSlwFvKRkMoqRUq2a1LYgUM9ezdg1hXIdDz2ue46S5ZNS8YSwSrGEr4gl595+z49
3GrsAWX0QxyGNAibNh3FN0vhNwtJ+KeF/U/knW1XvwnP/7BbHPG5YhECK0iPk0IFcFVjk+r7Pcna
24xtY/bpSzZDuZwUVwFJeaMBEP1hP4ZVW0j3Qu5a8AsC/AULBM24hhiWt7aBXvVP5BoFpd0fFTt1
mAgkDdJztsx+dzZnPKODDZjPoZa4xFPnZeQdUTiWdPrkY0Id8UtBQ30b2o/ngu23ihz83ZV9Eu/e
I1JkKIPh15o95nhWtXVDeTFZwaRzhKTrO4aQpeO331Ha69IgqHcS7VzBYMpRJ6ToJ/rdPTIy1HEy
xb8E5V58Wjl5cbDJBQBhI0cZ9+vYCQDOzkYpEiiS15/CFhlte7sD8kfrpqFDzFjP3jvmV+0Xi4ex
rIS5H+xpVE2xdGkKWiellB3+QzmWYQ7M8IO43sV93k2MtaTevYqJlr+amlys5gkzln4/WI8Iqqf7
TuPXRPY/LhivI+BZah/GKjR66HBk1avXdi7B53r3Qlix+naCNZH2+3yhPrCN6Ntx8p3H2s1UelPs
rI+5wAO8bgAfSK7Y/XGkoABrYjcKyzz78YsnPBPsUFywdlY5c1yOpNwhqhabBQ8zMCyX8JTIRo9x
kQuJsST+j8q+n75xJm85JHN+ppTbkETZ36PZd6/i4pi7Ek10MlKu50/Hxiv9F7ah6Bz39jDV4wyU
RXllQd7Y5WUhZe39bkV37UQL3MfRvN9jxgyt8pwUd9cav6L+kbM1lpSqjDkKxMhLOLq2CrRW2qdR
+E94YYU1j8lJipes6CultrZc7rCvyPXHlrRxK3HoB/cyQJCetfRwShgP6hqtpBHpuJFsTlulJuGR
wFH6/6onhReYU+NSTLRDXcW0bzpU392pVBVTEAFyR4Z6eSUBFakm52i/e/pwTvMN68s4jQ/io6Rs
hQ5V8MmyhKL/u4nawRtBsO/Omz+/n1wdmJ4X9rkXI/2xJarA+MB6OUltiYlDJkd0HK0SxySA3bnm
uSsr+U8F4+wbid9WiJHR2C6pD1YBpz9coGxB4s3TUMJM0ilGtaMExDCj/O98+FMk6o05fJWTdA9N
gUmmCyIcbgG6w/R+jc9XXdOM/sbn3THgWjBmaA47M/dGi7Kba0f4+x4bUCFlJQ4MpiFeB41Mv7HJ
f65R06nYLcq5ozJL31Iif8cFisnlWLrtrqj4TapBqTmT8GK29EDf4akSIvHX81ZByoWwgDrefMNs
olzHySsYJjN4ClKqoMWSefGTDpDOHs4NVRJvWY90Qa1dwLaQb9nN8nBKFwVSY625thyadEq1XEbh
a0l+RFgCb2hPffsGOGUWqyfh3jUdyN4tYg+aJYX74+Q4iit6IAZP7IeIPBe5eScDprO3VZez7GY8
1EVmu/adiqulIhmISFGzvKxgvvHoe+21BjCJj+mmwfeV0aCkpfXoqo4rrBM+tujZ3/Kw3W4GApdG
Ik4Vvw8vFVfkXHbibUdSM5vr1tFugqEghTNxnoAy5bnO3mwDNeTyM7pTn6f7ZRuvV4md/jfkRVvd
e70qE3VbkqYWD5H6+52mn6v+bpPzISOjxm7TJYYWTl6eGbAeVqTBEJHbR0XdFHLYeaPqoOgHvDHc
p/2kzJ9rrB5rfhTUFcvHxH05dR0nYUxwALq58nKP6yuXrjjaCDUS17/+JTSXXXJXRhA/E1EDz0KK
pMVHBk/Z26Q/1YMVHNTgzc3M40Ptl3Uiiha7ENSajCmdjyA75VhQvp1ubyfKQNUfnXwraM8SbbM6
gbrUkij8OipbREUvr9Recl1pETlSJtfVOA8oeqQqkgedREjdgw928PqaGormL+NFOqd5vjtWbtwG
gONiwqs3R/hciJM24W34IxAIPIqRHsVPaDbA5Aj6dNpDCxAGqgtJG6IrteohYLQZNJub+jhZsz1I
P/GNjZJGp5/T+n2zXmU7qs2K0dNhjGoQQJxCb0X862D9givByEpGD+For1Cr/JUXKj6Gtqb+iseU
/4KQ7S/dAtSBUNWk04CWsCU9xqxhdEvW6gkTHYzFGe8KeliF3LfIKBX+XquwYTltU1237SkDooI7
W8jz6Sc1dAy7DjKHFWzvml/RG4NYQn8e6Qy+F31mmSvWpo2s3XxGwJTHkOyLf/3ueOo+/AwMTCO8
oreHAVPCEUcm/Ua9aEvOvV2+EsHcgyiFtJsPfKp8FK/xp1xGh8VpIstJ1I7P4EzGuORH5aXzhsVd
TL0+aJ5rHC51kI4ezNbxAj419CSuRFryjXoGO9N/4z52XswSK7rvOy0YxFnt4MilCnjPpO61ZjcQ
GPmYFAjX5IiZyIYdfM7v/SsvjSVO0hQNmkWbAliWMwSygVuW5CG21lQsv24rmEztb9ZZrC7PtEut
QB2119DoCeJ/5FkiM95N7/7BuwTNC82KiBgiojIbyBNWPoohK6j2a9Nld59xCMKDyJcsJTbXoO4T
jYyYYteAArNMokEfWFKWK4PJtjOEMgu68v3TqZeA7n2C31/NA2QSpo6+Ym+TwYInFN53m5iBXyPo
Xs2mJL/PTQW9zmLuiYldPDXxjvsSUW8hbGuhBfcp7pOLP9R/e0O/aEpPBkltJeFWWH9G4kB5tMyg
/aWpvpQLF6KCVBWXroWNej5LduyFS+yU0IyHApH4sC58hKurKMkTLBKXajTNOwdvnOPVYdr4acpo
nRhJ5uZghCb6gDcUp5bRpwTKYieQM76ic0IisrwPEFXnZaLwSQ3wgPsX7+7D/Ek9Yy782lIffCpR
dk6xINLiBcG/468vJvdduk9ro+kuDclTu8EeasBsLqd72dE29hCEaatCps4HBREX6CsWi0Eifapi
kLbci1qX68QLgc5Eg0FTKg92XeMtJUHd/209iiQtVwJ7PulSwPw/inshBFRlMflXhHeINS6QtUcT
JWb8X9ac6CJlRgyUQJmySy8VpjQDDgIPldTOo/TYDRexzxgf3WWNVHgWyuq1OFrURo2vpOan5cXI
Sn8C5fQd4ZYZ60vdg5W1Hso73Gb9IV/tqxekwFJIInn7khle3IWaxFgAsQEFnyqTIojUWLLAZJO3
0DtrwRRhgRGHwUD9YgZX8kXfVXs8iMZF0xniYfJw8fecWuCL4vBmJ9r40iel44u4dia8CuzM3Amj
6OU5kTwWmc8P2qMP/GVmAnAp0MI1Q974guk/Q0W4Hha/9eX3RTGAJXJTpGvxcsfVPgQQFCRV6wo+
NUd2mUNizMnGpvMLU5nlVj5p6p3ef+J69ugTZMWCNWHBzsSAq2hjXAsWR7SHRWULq306tKAFey/R
gC/kMwIzlao2ySLNI7vPf/5FIdXPb0Qq969MSoBdpe8Ir6+ixlCyTVx/4OPMzVzqdhDClK1eX2OI
kdvhjGr38kjEnNFfVD1cdF0XrR9V/ql2VpKLPcwZpUIsUtHh5RYaIg9+UOUvlu4rc8yBvs2n0c/F
O47VkOahA2LMd3Gy64Cd4jBpuPethIPuP8X+5mY8084fpBZdWV8hniXeQ2/iu9VU9Ko6BeumnFGV
doltsh+MMq195/0MFjZjDq4I/u+Nloldp/MiVj/UfC0+nmPRkJPbsdTaUfLVsMHOa+SV5dlJXUel
UoPdrZJZVyXjA4osgEI6funjP6x4fIxFyJk0PaXKmJ+14FU5xHEe58cjDvDALzQZ1l098ESu+41t
DXJyB22Xx/vWuui7R1mivr2Azp2mjtkz4AuPtRJRszfT6MqbuBW4/Pt3LsHro0H/KCA5ViHZYZM4
Ndw/GFSrwQbWdWUGNjIjIJSZmQfTwfH+1s+Wq+Fz+rlQvn/9a3Hdys1ZM+WTX0b+Q6M8Q9a9VweH
1meW2zpJQ8XKlXPN1EBzAflpzMWtmsN41duhGQ7fwR2a0w+RHOD6nS4r5LK9xiSVn5kbxDbdLRrh
NIBqhZhhbGQpwzNuOVeDWlUslf6qYEIK5sdSj0EK4FJ7G+SzJ1HMT2QMdIysPFsTfZBGUK4kBugu
mvylaEBJCU2lBlet84RHpo3CH8C78ieR377+znGtV9twDZ7uTsTz86gbCtnUbfbLw9IfUOmKtbSX
F+OVXsqk1RK0LamteCu7gnc64W6pYIi0gyT/KQviSbdKkpyxHtG+Sc+phJ2xpAgDYHx8ZMZRlHWg
E3wIWnzTeLx9AwhwxPOshFideOFc5WryFafBLqfH3IXWvryv5f9MZEhqnpLdmvcD0OERnOOE2kMf
3WzHQfkwD7T+F9wdD+k6RaJ0G+L6zI8jban4/tx8SFnyrY/HK3rVY4HMlrJrf1YHfkdhWjPQqxVk
jD1bSO2k/1ADUGhTqXDMHdTyjib8U55jU24uoc3Odkepqy0P8qtEaif8oMwljUP9L/bfetSr24rF
Vr3Ud0d13X02yKKIAuWfKMoNd6H+xUrjXU1Mwdx/POjkdvySbNcY85ZWgkDc17h2y/W98w80C/ah
vbC1V89uld5roWMAOZ/X27yRWRI+dTf0QA1y2Fa1KyTdLrWkdjOP+G96sAixRWPLhSLjH/1pCzWA
XaNzqRC3z0AmDm1YtIv/Sye+5vJjnw4MOUFFS4xbGDueG1kLLBy7TYXEJQBnnGnI0l3bLoQRgHCY
2DfBfqitJ1k2Uuxwwx/Xe1Mcu8tbRPstpFr19WwWo71W4vF0qCLXbieHNhg4sf9h8CmuaKlv6I87
V/1IWdNTUXBj1Fxl2XZ+v7J+cY2P+hhUmgwOUiDKdIZGMaPv4jQJMyFGRLlgqCmrA/SjEI4+hO94
djiwrKhmeEsXN4yjFaCILr3tPmn+frImsiYA52krwx7amJwCtjdVlBnD4zHlZdeBAAXH1ZSVGpGo
iOJs3gjM/Uttbc4WP63qdpMGdZfK33NGMbseCSvlaIItVk50d50y+Gn4aQmxy0oPcN24zoYGM4kv
yLoqqcg8MiyfY66YZAa8oMFxuqafdpjIVtU53dIGXahpdwylGNgITdWX/c5z3Ev8ZSvukbWmtSCK
I5ZqR2cUDVV4smMPFqOWAXf6DiQdSTN+3nVl5So6ZQENdVD6W5LmFnKe2MYoE4mVncD8lR5nfjOz
sMnPvD03Gs1wqBwHa/D77xPdDx8+znz90sJi9d+bdPxCrKa37apA8X+2NuwJOStYOlX7RR92WG78
VvV6nZ8ZCHSVRySWIVQxZH6XM1JUnlpOxQTSetHmxrLdvPvxhvwJ+zrRI8D3fPmLnUcC3soWFZVS
KqCxTvATRe9hrBXn/FZS/ij9wUwJWrHauIhxMBP2YdJpX5kTLTPNS7Z3Nt/lgDd/c7tPS3bd7uQk
6gUkofyJangv2/1S+X8zUgRUHLn2NvGN3YZwohBq5y2ZXJS3uhC0uvd2K+RixsSgkXX7oUDkWFtW
6arWPQ/CEwIOmwPXKICXduNULZiUT4wGFwqjs7FpiNkU3Hr1salrJ9cWFJWF/JykLa3xHzenPCeJ
LeiyrPUwLLivIbRrY5I5psx4FoELvij6qYXtEBtzw3xZqre0UyfoQgm013sOvoorahp5gqKH1EgE
ALCQOohmqzATNIJ/965rHLCOhtBJeoy8s8R6KlGM/D+k5nPoMuoclFJi4xgUawCvF65fbInSG+7X
0w8/UzLJ9j9WVB34pPOdoeFfBGKsAwrae08X3bmpu/DQz9xAU5btezYsocJ4Wcw/5Cc+8IjnzQ0M
fT7Ir3AiMCqIGgsmZX2TcXE0pVhclL4CQEN1W6xtmMmtPlaOwD30vu8VArEQbG6TscmKY/UxYgEz
tr2ksHOm7SVc1RrUulxukVyRU1YeDJ+y3Zabn1gcpzKLuMpOEDkz1OA6Us+rSQ2zNOw8Rr/Lcgmv
HRWXFOtfMy8uZi7Og0fEv8qBhNIBYy2TCz5oUDyuWvPrwJNfzGfub8QqQhEclYL2lahqoSW+38Dw
WzqztNFzYOymRa11XORb2cBzlGoSXbBCYdWrJWGp+94GiOeu0CnV3qr/ZxQv7Gpr0lMFhrPm3uJ4
JvRlOfHPFV+VhvPiNheXHoUQd5gaq6b8fKQCOmbovcnnbPBe+IzcmpdorZO5IwWTlkSxCDpE9CdD
A9Yfn843fCZKvCz2vSuwfws2guQtoL5Re2PBAE6cPA3dNX+1i2U8Bib9Fvqs83QbZk66xofxBEsC
R0Haj//kri66UP1BTnpSGJp34YQ3CrQhtfLgX5yPI0h7D8Je4A3GrRYnc/R/1Rqx2tBo65wQNozB
ioOTw8plhKRw/Ayh4AvEOngG4VZi2rQymERqegMJNz97o9arw53EKwnpDPB6o9vcylQOcZFoRdsO
it9PPiiqfQW/bCJEMc0xWHO0ycvRq0qHHu//iHCEM0An6kAy4yosMvOz6D6yGAHS3uieSutVjAdP
mjCtkOUgyQ2p67GRed0K5D/pd0TtMCCkSgTNTV4kZkscgoEXvAq2yR2p0ElXgZ7FxTFmODPV+ExG
MvKiiF1og+MQWL/yiLvjdGgrI3j1r3nd4kgqZaiiFSxznSql0Pshh+Kgi8mGZQ6zU9G8gmsvI/3u
qDpLisSZh+qcbmEPI70xDfNb/hg6yNVJkBVUjaXY4ITJwCvkELjrLY9gynFqxUCPVgXciMmLCoIS
WA469xmhJPC8sdw2FBrz0kP8qFw0SEaCQYJ8gEx41JIR00meO6R73yXhHXFvrVo2N3PM+ESVnsz5
3eeu1/XNMql1K6ZytAApuG7f//XvfjnHiV+qfe8CiJN4qY1boZUbnz4LILFxZsEWUsXfbzoxhjPW
FCvkaJ/uof5Htzx7LMCsGiKtTb7AKbLA+yuSR3l78FsUbpz6jFssFGgz7WS6Li8UCr+Q8o6l2dn8
lnFJl5xJE7/G1XdW5SwTZSEVayvUthIzL6KT5v8E6gJszo+anxvIJsT+e+t9I6SO+O+DZ6BGwsYa
jsZLoRDkX86elnRvaREsS2ua34tXhIM6wo9ec9Tw2ydUpeSeD5Z33FdfkjDW2rYG4h8ijsT6K5vt
UIyjkUgmH9zDAHG7SFDdMz43D7J3jZOi9IkuFkhcpD3WaijIeisp58X2ioY0iFSXIxDxGNFAP0k5
IU1fG25dsZBp2crQB23DSN8adH2qMWt+NfHOCBrtBXi/znL7fYvjXmWMPniaKyn1zYODiSsfk4Lm
+BSbgGHheOnMftHX5SlxE2E+uZxU5vuDyU0a0WjK9KOOqvFNd1H8Vxtj0p3stKX+jDYbEPVxHHn7
ZsQdoYxkMWn2/W06tIEot3/N6FfKZtnQwI7ROYgqDUCl4ywcdtXhFMRux92NAOhvft4BNOPYee9T
aAeeg82fK3/sdyHkyPI7naQ3YnsqD0Nl5myPnvoJVQSOY6I8pvtKNRPR785PtIjvczE8Z3Ewt+0T
/zot6cwKRq2u0mhpEiVR7g/jOV9WnBGCyr/nOdPxEwH2PEvcFq9wczCWWxpekmn2cwjuHbchu0k2
Idbn6EpG4v+8OMin+w3Odsnv4mQxzYdigQ2JAHNBXHW09ivwWW9iRDypZbxcSCAKHUAUiCyD6FRT
OpD0JmPtNXOvYEOi5yXkPPObbRplumkCmuh/27ZalnaP+jhjpy/4+ywkSQLLXSEqPVwVUdJyBnba
1eGlEW6JaBvTyezTYxGQzArgKKcGp/oxrMIlXOKsTTczfA7Pnw4fmd0kvN3+r3QPrair8cZKleJ4
78yk6skpEkYDZZALdVOJHsPQwF9yA5yDFiQc7Ywh7oZZZ+28uyGUrKB1JJKMBvXB2HyTDPNl07uG
7RikdIVWSbleQ1LYrp+4bnWiggK2h6FNsTZJoiF/vA5SxWj+059Sg6k57GNkQ2MpjB26b6bTzP4x
EvU/vawL0gDoBESYlSbyhfZf4FGW0E82+b+SVMtlnNRFGx2xeWOTvI1ByV891wxDcQt+edGMqm0Y
OrAS6aEy7bfMiHMyX85N5I0vQntK2ge1Do/+exJJc+AM91tHxYOtx0W0XpBtGzpa6B/mJqq7Hqs3
6UFq52rZeNb0hdEcZ85ylV4e3SryuHAp8gsnpXLxEGNJ3OQpBaZl9Ei3T4B12HVqzELf4SSLI49o
t8aPU/hGRLCnJXll7h9voQZ6G3cf0vRSRF60euX3An09KhJGCE/rscYBA5nmu5v4sd16QE3/m9uc
S585TR3TR6gAvOMYDUzi2hQ8KS3yUbDmjRxvsgOLGx+wztSDxCa2lImitjLTLYxYaHIHdjLQ85yb
fxBIVmpYJ7C9Wr8euZ7psCUoRoxKtZgmzThQd0sBAc/qIJtoIBz0RH2oQQFj3SIAAuZmi2c8ncCq
cBgAbDqRS918m2/owZQ3PxBJc/PNjnqjhhTYcs34tyAptf/Cb76+f7Lv/TmfJctgPMltT9Fe95um
SjQcsjtPfAV7yNV7hJcd8XGJzmz5fr9tPqudch5AEugDtM9ab4bxYyJzuCFuj/B1V4xZmk2/f4qv
hjPFaWDu3HOJ3np/UCBFrGGbC/3/tw7McaSxmnxADDsHG/wHcTZPnljBj8ed9/D+BMNlYjRUdTKn
kvA28hEJcKQpeSz/DASAFcd9O+W4cGJcqmq24mGSepzOIGWOguR0Q/BSgjaH1UjE6s46c8lVr3fZ
OJVeXlHBV7gd04Bmy22M9VZ7pwjOxkTnNzFbsgzlgKUAqH/WzOunUteGgFbkZT4bMSvcvjnwCHXa
AvNp2HsKaBhX38Zes+VYJ3J8qDK6JAx1g7IIN+yD+xDr8sChvPuV/+28yFmSdsZ5Q+wych4Mvwjq
cX7tIXu7GKM5ir0tEGOjS8ouPvUMtorGhg79SuF8PM2MCRshXb1MWb5FL71v+9FKuHKJB6ut0o4Y
mSdIxm96ybIZlZPWVegMFoow0TVqAoEx7Uuu7mtQfnx3RPrHyosZlIKM/Q1me0ihHk9QJFjlemZ3
Rt7LmvYzC6fuiS8Q1rpAYar7Dg911T/YoNA+X0lmDxLbmM5hey/rkFzUgbys9jhzrvcR3xcwrBeF
EZWVTKJWRXpOmy1bdVj7KQtD89Nn0dry4F9mHvEukyUTUOjbd5ihf5m1fP9sCWSn6PcVv7bBSnIQ
TIVI1bd+zRotSN3sNWBBpmE5kdUzbRvPcRYm7RgbFVzYboNuqc96zivhzBTUL7hr5enfbBHtY8c8
IyreMVBBb/vRZ4wiR4BjkWsxFa5hNpookbLyEEFyjdbB+rhQ2qH9RcVw2F+Q7Xi+fb8eF1ExLVCz
48qPMuRcGgBKsQfvTq6q3UGdtJwbVJR37i2FeCYKWJj1YMuaswn/e2YQoVnNqJ1N+cgvuek57unX
rmzYNOsoitNvO1PoyuVkpyDRGVFDP3A6Isw3BgplF//FThNSMu9qkV/WFD6E/0jDwc6fNG3hoisu
lu3JMwDzWs9zB+AKjEC9d1j/W38Qtg7BUDTRIycIO+dyx3XTdpypeKZ97qeDqwskO3UufxhmxmHV
7M+JJU9aaz386mcI4Qy03c4WmhqSvUCk9tCkovlQkG3sHyc8MOHzwKdE4ltdST6H7wn6Duz730V/
b9BKD90ThEYDogHN6vJTxgNmmUggcFwl5xfU4/pQtBe0Mg/D1fcEtrU2sMDbPD28r3O1AYnQZg3V
bsLJej22Epe7MbQo+v0my+3Mz7Alv3jrWRKa0fuVbVCX6BIruHqyCCQF2CBzkWZxh2X+A9uQ4wFu
A4yA+EHpK+Uy/8Pb5OpOF0c7RSHduIEqYSzPue3B3revgFj62X+i1P+JJWw8nP7N4BPsRPv5qMOi
LVi2K7hAm7338yjiFMmjcbL5p3FNkH9QvHVvwRYlHH62XKPXdF1JKNrcOndG0OqEeHFaiRQD5eUa
3Ne2hzKoPEBqErGQSjPHyOXOoZQsP8z+3t7DFlZ/94tH1okaJb9JShPVwyUYAqvvg6oW+qBAUt+G
qzrtqza+NTB6ZPvdglxHqhKJ4hq7cJDazIEgTE03E51RMOmg2ItY/Kd1UpuTlz09RkqMjc+P2Qn6
yHlECCxK1jUIOHznFMiGNcHATIDjXQhb4EgGdBt6Fl0qlp9zi933fSGF2VvjJDzn86DfFKyLaxx5
VasNOJ+P4iPeS1pnIzzwXeTphqfDokfkorD8mFBTAbBs/hLu3Ts9kvnT70sR6w2yJwCUnSJw9qK6
2LwD1V97FfLUMXXdBfgNXHH6HFAMOcasBVakMsSrlUT/hs9aW6SOMvpQkvCT0aw2VGeRgRg1KyfT
y+ZYsLeYrqlYAjoyu406QHWMxrf00Y5Ghyp7rQWPobMLMo76RYLmjJMmnY5hbFirLpqgFwzg1lwy
75dJqdbiNbfsZWJQwuES1eufUbWna5R4OV/Rs9reV1zzGrZCAhefBk5N1MiU5IfqFh1Ba7Lax//H
W3DI7oLIC8imZqSy9ojvjt5yD27q0zT9nWxGeaFL7Pq0vH/ZCWiJ7UT0ujO4+24kKkAUHcld7eNP
NRhrwZ2e2ymCFhajkB8CjPpYwj2R8B10e+zaSPp4ZtOE6MG549zgxHlBJu+UTOHstQ36yPSz0Yb/
1CaEMStIyVGxnNe44xGnKbgQDd0lSpxZBHXTcGSsPU9sw2yBAN0ACTf7t4g5F9oDCkc1thjl58M+
qO1qhcu0KDZUq7/DVhjidIkI5OiCZDkR/nb6lbauAvGD4jMGtJ4PD+DngMZjdHdnyBeY+jJMKiEK
DCG9KCUXSLJH+DlHNCtMZ89lPw5dSNRKSC5yv8j74Mn5D5xG0QW/urAnyeYiASacyd/WM9agAqio
zaSAzf6hV6IsauLgqHU8xVgos+Jz9ewvtFnAem00LrFwf82SuVTSkFVlX5DkAO+uwzQD2kO00rds
vLHTsM2V8LRfraEc6j6vq+2yDb8uUhmhWZ/0VKKbvay35tFDZOklPraF5udq31DX8+CG5TdaTc2c
ITnkNsjKoCebTDRpYdtyS5hXrfjFEqoDTRcP73szrfgFuf7/UhYz3Ye4al+hVPlxumgEjsVm0+5N
ywyDapp13A4jh18t4//M3wwBfjV+VEsspXdhwZHyfbS0tdPKaN6wfG7mk4//Wyka+twHP86ISobE
c9WyWVmmjQPjvA/7hweyboMZpCIKnQ2Z/iu3q/BrqNcSFC4m8fmsiyqYAoJ+NGECyIGCY6LDVRBp
JKyAiw7RSrPSp33cy+WSdFedo5RwQKgvv2JA1pqWA2lXIwhZ+DtoY4JisT+5KFC3dNMcfNUSP3fP
L5Ci9rOnd+HY+2k83Gcczf+nZjJ6LR4fMGOwNZweXsupBZX3vYTDA8HMkIl8sJ0Yrnv6uCaYN7Ri
2Ce3NXf0ijaSNwre1ZOO143BfbQuHRQnkCN2UbZWSFqRqKV4KqWLuEDTCH28T8T0cd5uvaNjGsnp
tHxkGWpiY3f15IkdaDxr6EE2wh++sQOjOfnC4IdFMywF11MMI/pbOeRaPylc/XJT3NN5DV899eIG
5QN7wNjLSBKRsej9KNMxgYCiaeIaK2nQHCkZe6t/YPOzBdM+ANZLHHbgxj51iCkDB8LxOozYSjf5
P+Vx6F//4dSA13byN96afQ0NktfiNXZEPVXSDYVXQjDoReTOH43lndQo7L3yW2n7UBxg062nOtpl
ZyqGLNrcJ9Ao3jvv0AdtYt7HX/mK4wK7uQUneR9eAjTZLaGLbqcMbTZy6hOC39FC+DO3fOQUx4NM
/WjgvVe6RcwG3ufsPH+FZtE3j5hqAgQ/UEPMa2Re2Ht/XUhkK4c/56pquQsEWixRsVeJ9IdOI5J3
SPTgtA8FHDP4ODr/UM/TenfWwRmn9+/3HpAgVpzNlMVMgdMxMD1QEtnkGnXOXYmON4ujv+V4rWKo
19/4sZyqS56BjcwMKRgSFjkrB+OUXijfeN4bnyU8PTQh9BwHXW2u8gDSTlzQrKaAyhGtbV5ubdL9
jpbOt4T1crGK9+8IZib78lpTwGFZGAlEcfx6GDtX/3OV7xyKHFoyRt9l1ZoqgN2Md3JBtHLQ7X2K
L69vIbyWICBaa0UVCgoSHTcuUIi/TxITcElR/+MUtn0EmMODl4OcZATEEtQPMsFuhRibF90oSIXY
Jq98PF+FTJALgzrKG9ktlN0WxLTkWiEeSHvbNwuHVjjbG/wc1mBotBwwuoN/0/+e85qmMkwvf9pt
R/wQ998lAbQ4bcrfrbUqOHl2ACnN/DrkfEvgDU46O8mkpW2XDgvv9xMp7a9eyvkJOiRKPdoKn/Da
1yYIYlsNxHWk0QJN3c1YZVUoicjmUU+yJH6Qvyi2/+uHGBPdwOptiowfxUCx5WXiDRoCQoWGCZXC
zhYK+zVf5ahyJ3qYZPb4gMI4x9gjZSdKnlx0GtoYcgohGELE0hH22PPMFdsKoQC5b6s6i/VOtsjI
MNFkGV/IknsdLxV6KsyVBeCIhz/Wf6/3Vh3F7N8lXvZk3C73wTQ+Mr9ERVwaDEQea3enNISFh+v9
OCN1J0k9j19cDm+S9bMsRRzGNwLPUS5TShVFKa02qLK6bn0b5K5ys0esy7lFwxDV1y0ZyLnuYyro
jf82dueKQtw74H8G/UamnKPurVW9SD6kiXpSeijGBwgThPieq98cQxXGaQfamPHoYtoyVnF0xcIv
l7Xk2vtsCN2OthKwI+qchlPTlXGu3e44TkPwQmuEnuJoeMvpCzIUCQ6i+sp+UfpmYM7ejYotQv1U
7PUT/z6wXCBun0SjNPtPQNggNjJqQc+T472V4OGJfzhVVXAg1URrt+1qKHjy7sXcO5WGfsipGB+H
rW1+QsA9PdYgmmyD8b7s1fJJeEiu0aUWk6lsja55oKZNeutWa5FsB+vZMQ33XyxwlZGy4qBuaTBF
7Iuiud4GtsGaqTcD34zl3XNh4OAVidDw95zKXh+XvUsx+uA2EzOIWIGysdu9NWERHfc9uubNjt4R
e8+R7HQFTwSbK8O0SnJLz7tMs0WeD6rCQwhDX6lLVyeWQ+Ndxc60TUH84Th9PIZ0CEQf7MP8Ela1
oPV+fByB4JiwrraCZNvKV+SPNHS4Hpya0OpGwHm3Aq0ZY155+8J+DWGiiwV1N/OMO6JsP6ZnwUpE
7Dsoxk6ybWiiG9O8Buq9Nx1yu/3pgXPUz+pmjbAfWHb6bc52X9pm0yHPYumBLsrsDBA9mAYon3/O
S715GSMD20C+wCGG/+/dIYL8BEm1hL0NnsPJsB+OE3v01yvWDKxGVd1otnoacKZvu907wm2ZcCod
wpZoLY90k4lxo3qJzrbOWSBfnExfqkvelk9PeHxLc7lFaqpvnlxYdn1kuWnmUi8OW4Po1Xhb1qYU
ALhjfFfN4/GFiD3tSB43Jk3IcxKVnQYQjZZjDr04xKy0fxkJTAOqOCjSCUfiK1ZehG3DzGpPCX/7
q3AeYdQD45qZ1q84wfKkMIKnz9TYjhBLriOLjmJd97sYp2yWVrEDsVtb4RwIQdxBvey9lhOLqyI9
9bwsBgNeNqp99/Y05OyW6CuVB3IFong1KfHRbrKXW0kb5HOIsERHLqR2GV2wV24+2Y5/VkZF6Wm0
EJHjRty/qUi0rZH0Qscv6f8mMo7INMt+PkRJEeQ4ATODfHCT3bp2Q2t1QBxFLAxAzPjKv32NxMyX
BQpOQXZXI+10MUrYzu0v6zWgxuVY32jRdFNLp0EDuzRPHizgzlwnZPs49yh4xvEzuGjT+vXkZ3cm
2RjYXUMz+U6aBu3p6BI5BTQa+rQu5EYQgf9qDx9RIF+d3DpJz3vfP7/IbAED0iSK/8XLkyTbmzeT
1kKRHOhBQTP3ML7zygSwYkovAOJXS6wHUWVhbjZrR7rPTHGaHwxyht07pCdrKIdoPIgsJ5JYo75M
lQPQi+pCvIQ6E9g+sL0VfOuZhkvEdfidROh3mEppgmDVf3caeHlYYm8ZYq+zYc+9ZpiBgqg/Dorc
DUl5KWqfrj6XDOtnUuv4z8ORMTrRgCVPF1fRKAwfFyaWbC0KCdazNVVz5xFjLI5P04GPYI24uwOg
5NpHYqdAiGV5Bk91Ljj9OLpc9fIutDPuWRL6X28tTKpqPb+J27ogdUoMmiydgYmJB9KAg3L+YOcB
3341iD6eG6d/dLIAaIuFBVrV/L0L2DttCDGqfdo2YLZtuMfCiim64aJ4Fhz4SxstkSsj0EooAZYE
UR+a8h4hkeZnqXe+gaEnjERaOq/6Dem44iKEHiIXBBdmYvy1RGLtRrpIcVfDVI8JSuU6Y+Q3nBpz
abRVMOeom/GoOezEWCWo1hCEYut8B8qoKWHvmVpGwUYX0zSFdHLsy6tgFBn6pPJVCWSb/VYryqCv
1lFEIbDTnL/NOqP3NfzCJmD7LYkWCZ+aJVr41BfhDgSCc0VglCwsDoCdmD/AANpoYigyjCI5CVPp
/9BQ2WhpKQdhJn7kNTA1Y2AoKCLrBLcKuUWV9H1zzjXwcKNN94py8wIJaR6kL28WwDv4T1URw50e
9omU2EJmwolVvcmbbc03PnATdOfLdC/a3iG8j/R9WNcTvuZGdv2rn3sNHgUr5L7kd3YMQkJxVZmR
T68n/W6XN/o0pfLIbFOF5WprKj+Dz6jO8KrhTA3pp+1t7dSMEA2qGD6DzpUXF5bNIi0gBnLxVKzs
TVaRiq/X+LMvvWQiQcMMtaXRj1eCUPm7YM384/jTJv5BWWgB6orDfTswXAskfy+brW0xK32Xt3tB
Gn/v2whK1om+Rlst+wgLpVmLeOC3alsNNzBNuwWfbc8iXWuUbzwb4yrgX8pV/zuo/79AS1muI/z3
phySR2zn/jHfZBt5FCaCKteWVL4w73Y0lIzxX/NH7ZPXmk5Jt/mBWuoNQQYcPhJ8E08BJ5HvWeHt
XgeSOZVO8WR/egEf6461lDEAvQ9Vh/mRr8kaAXZNjbKByvxUyk4i813hjquQgAquPsdkXpgYhk/j
b+HFIhYesLhE3NE5PbtLGmN2nbTLm21oiIiHhUmqXjhmVNqosyKhcOpS+YxXtsX+qRnG/Fug6lOy
vKxqnog2OatR+ruH5iKz/3KhXt9IPtS3wzTGaABOGxRY6gjYbtH0+2SuDtKmQqdK3eSEj4nSD2Vo
MsDjGq6AobIEAyfOssDKh15aurSoz19M+GNvEPQYOhAzYxomkPNEAX1Ymfeu9QCwzMX6b+/MEqKv
l6uWxSx8yPfPI0wpvyqUJAer0v54ZqM9dLNS0/DhR/C44Km6JDfQdxZG8z7eL7sChwKQEH7EEVHA
Zb35VH6EGUIlnvHEkBvGg0NasfcF1f2BqAu+YeRhWMoZBs+Kv26eWtSCrtglY0r9CqPrMTlzCoAv
gB5UrrEnJAzgTrUENsSBDltoNEq8xgujN1bpxh64KSEmMqL2QMDJE6wwcyavlstNA/mdyNPG4QR/
yPBWKHWZDAofuSOULAS1PShM0VsT5QyQGTEk+lXhCuT2KYLPVzOjUhERy8qklYPUKQ4/GNTH/+oG
ISEMRXQmamdA2Dn9CJbaBFfBDmrt0ubFRJaY3mQJgXj1DEOxjdnHiwP/vJr4qyXrm5QZ9VBmezxW
TKST1YezywWGRVI3zwkjzfJ329ZaVd/GlW3gN8h/bdmifd5wWRUOs4DVJNlniSSR5n2fUBnJHo9B
s6i4jZPMnRdYpdIFo/mAoD5bydCAhRWBvymwABnEbfq7dJckTGGfm0rsktDNeq2aTFv2MjmbgsFZ
6g96sWm/I1KT5fmNq6KPrMLaFXLvWKf1rjyKrHD8dD+hvSiDDY3pZAvrdmRCBwzhT7yrTA4JT2mH
Qk5FZSQtAHDE6a/XAytUkvAxaUQAZJDnpsZwz/mKYccyEl8rQ30zP2mWYarF8RjAigyb9GTotNvc
faHzkhA7lSBX9E9wDMSjxU1Ys5hop1QL5cnOz2UqyNBrgJQBCqRaREGK1KptHvlbz2xAKX3ao1iM
hjFS24sr0xeitL8Hq5AoifSf/pqIlww6xHBZEjf3oepwbitlLeB+W2Fe3FtUp5Oo3LaE0i2wSTS3
CgX1qI4gXKzMxX8WSW9cdrQdI3RwW8lUJ+HMkQSvAB8afV4rR6Uz+6oyhOlxSnnXiLaLGVbIVNrB
M1v9bycsqfCIOPBN4D9wFryEoj0j3q7mLkhBEohvmiwv1qQOZuZonudI9AsVUIMtqHHtY0bS7ab7
SeAbgbtRE76UMGO+KIebu1j5I7YR2oeKxYS3UL0CDORv8QRONr+Ws65RYd3yN2Kq1oyneQ/DRgBN
jjaRVXsiEC3ez3Dwuif/Qwk+Ysuf4/bs590jo6s6/KJXr4upSYyxRBRaYyz0ZA2cm3n2Tsd+wtuE
R01EAdgr3nfHosz+kjGWQdo7gLKHmCkozS8KlpOiDz4p49LTTMaTkfRb689YmfN7dFfuBUyhKHSl
hYIQPlv4aVuHjlARkTPdWDtkV61EVXZUTX1lOfEQ9gpWMf/FQ2/Ojw5i7uLYlwuLid/5ETK7yndw
Zp2aOlR4Fr/IZdE/OWWO0h54VubavPhdzm4FGipfh45w1fu2px5HAW+4YlerR8A6OFluuLdMWnY8
uA+o1gdpSkRI4Cn78pMn/KJ5vuO/7P6J7h2wKrlqgVoFcxtjadhog5Lvwr0J1EiLZs0nbYa6dVHN
iTkT6s7KoC4WH3DZ8X3vOSo1qT5Cf8sXbAiInbedw1Dmxx/ExqDqUWGsY5KCWeMKghBxGTq6cDA+
/MXKTX157xFGl+9pFxOdoWwfw0eWECK+Q+Uc93VjArwBjcwp229O0Ta/+sEzbFuKMDfojVC20C+S
98M8NRxxSgUObH9AcdNPKBULJVeEkI+fxJvMWKiPE2AJHM9oVU9aym3ZTvBS3CHHkp+RiLlMWM/Q
OA3YIx3H18+QuskmamKteDSRP6bm21INu/z5+69jOLM6OxPSdVvem1Y0U5SyFkxQoZz0wZ6Zr2f4
rzWcW0Jlug/vvQKHwXjSm+H6fg4ZBfwg0EIpTUilgm8cWauW1xIJsE940xaB+r6KL2zy5XqvOxgW
0YSmK4pLQ/9jzhTaiIAh1DBL0jRzZIJlV9K08XLxEe+54g4Xn06fi0+9kEN8qjI1wWj9svI3Z/YG
6vo8dWNTGYZ8NijiNPASgUfU0l1Qtqi5HRXGFesi5nvzPLJ7OR9E5mSM+Og8e6PdUbw2fGl2btnB
YQ1DdemoDlIoZOHd3G7Rc1FQy3eNALrng6U6ZRLSs2LUJp6jaOeLz+QMlCsQdWD8O1+6RTXmLil5
FBUGKy0eJaxyLddjOD+76zUKY4vatuzpbDGWj5hCYfal1dKej57/Bfpl9WBRkTkgN1XdpdPCmwat
u6gj6JMYga/9j2wbl9zVUV88zn5utf5KBnSLEHUU30HbWcZluWnTMFifBAFPgDiiGAFBJLNQcPhD
bZOsdzPXUUSu6bwfQWHdGn+f6vEVsfiWMILJGOWcSbGaQof8cT9Coglak61ydDmKTT0br8esfRHf
sxL3FOGTjIYkyDm10b/L7bhw3DxLOrcHIQGD8/qMV7SKMveL/MO5uLqoml+fsD2wBCoxphrdTg6N
/MGiU8CkyyibH0eRDBdivWiBEmpykYnBQOxCGfK+0FGqjhmKUaX29M7/6nsGK1jj2bx2w2BuDj9o
F9DkHwhMcqE3HV/wXx2LBKLRRHCsqt7rjXAnkQQMxbKuCeSYE6BSiDXiOB56GgP54mzmXvHuDE+9
2ySbWmoL+q8I5cYSAfUeeNEUhpo6NB8e2SjcAAkSavyM9snGVyCgMdhfg3BpYLVKCQ5J1cuAvxfS
rLHv0z++CbHRbtiUqoRAHcpw9sQLcC4VqXPzARlMFSRj23ekm+bYtMsrTiH7XrL+OOtMiHVUV5oi
41MuZjTRTnNqX3HTVdh0tFWrQW7L7BthhsHdNownCJ10FXEEwsujuu3Jx4nBBDtm56kqFzzTXpQ7
HmYUXDvDAmyryUPJGCrsmPVZPVbZLM/Vf/dBhAb+hvPc66b4RcW70KoAj2cOTiKri2S7NA+bA37f
mOEj4aMJ8BocD/9Z8odl56ksD9mullEenl5BQdGNFVu0UDOWtEoHTRChw5wTDtzRLWbysb2uarZ/
NI7txO2Qffg+tgZkcqTTtew+qGRg5rI9951SgK6MfpNz01FYvm9PlNEDxeSl1+QvvWKKMUVHvvJV
wlS8o5OLwiXmfEajb+pykIsfLITTYq61Y86G6A5fqFETCdDjR07SJWD+etrMLJ4pcp5PQfNJ3e7R
Zvc1z3Vh+m4ql3jVVW/g6LqmeS522xJ3RrOIkvbXZ386jK39u7QJCxxL/bTkUu7pyNFjn2uHY99w
RCnkAJeE3U2q6hAyqBKg8dQOzyFQu1tie0eIiMCtZuue4erfIzpW347L6Rke1gF1lB/idMp5XMR5
YAnb80ChktzwUJJRkUc5C/SbVI8OoWyQWjcVZDfTNXV7f8xScuuaMi3lx2jhl3PSjJRU5kcjDbX8
DX1+fmOfjNbIj5i0Qg+SNcJJ0XlavCtzB7xuk1mLez5erT3lZXuH2DG3W/GlKktRTmQ39eFtpOdw
/DrzuKip64jg0G7kI3LIbqF5W04jFIWc3FSMYrejUkkeU+oTobjhQy7ROln6+rdK98S+bzWSGoIq
DKyUgu7qSFh4jHOGE9/bRx7NYkV+OvgGvDi+nZMgd94pSZFJ/9t6dSO+uCtU/v/h1V5LgVmJz2bs
qhe5HkxrlzSurHAHWeW0jEQoUCZKQlZFtSl4XDOBLdXPWsrP/vs4iahqNZWMNmHSZyN9qKoJQQCk
MPn5MZwchZl+qgGH1NWA53I5p6bUB7oY/sehWrJh5xOHz++plkXnJWhoyHGXiDRfj9MTGWgSZNS8
FDFBudSdqVhsiA0ErErGSVlCPCozZJoB+YxOK66ty/feeEyUVNKVW7sJ4dWrMr9v+IA6wHyd0VBF
E4TAhvcn+zX32v5LA5aOQY1gZRY+9eXbwfNGWD6EMeb64udQiHloJj70kvDQVc33dKWIZn18r3/A
nDJepLsAT5hdLH8Dnaotu/h80FfHNT0aOiu9QmydyZiFRDRgpB8d2tqRrRnTUPPeAD6uODscNYEy
1ImQKabRV59wA0k8edG3LKUnK6f+Sm8BuTC8Tr9Yrs1s9M0Sb5dmms7Q5TqCd4yHdmD7ja3ZdETU
0HWYyoSntZonk5tTgkmzmX7oln0POJLwQb4keQZsuYFw/O21hhPbg4USZTYIAgzjDLtEU3jLCyzP
IXonuId5YlP0ayALNiWnJVilDxQ5vUa+VxcpRQ1wZTeQyWNdCfoCsql51Yk1lXBn4xtqy2K1oK+0
SfEzfDpeK56D1Oq0VKFFnZ90WJsFb9VQWqP6Svq2Uatc389lLthhen3U+tcjmW6zl5z4q5PxBuia
qwC1ajKWvIBXS3wyWBtlJUTHpi/7zAlApOC+yTZQpahFwBhpt1rDj+bhITUxGAeCl7NDS2uILthc
J5FW9qVI6e1vH5KyLcN2rwkUWe7kR+khR9zncHiGOUKLothHqhNmzkCx/8fJeULIQO70eHF3+eFX
/RmVISHwYT/6K0W3ByAl5CBvXDFB2ed69cGJ/qyDQLcuIP8yZoN4+PM+33vuntP4/e+WkOH24luv
QC7NlTE4LN6hdqU7ew2q5CPXOYe3K7XjNphDmycLc0wVVdfGVmFfKuLg58cODutA3NhHRpuoeqPO
GPB4InAPpBHfh3ptiufZNxHxxP3mjMthqpU2hmHVwt6g6Kjp1P+V5Hj0DVEdnvMRMSXHGP7Zyi6c
EZZwSFxO6vdyLWbxCeVffpoY0UTj4W6CrlKEcPqKsohU1JcFrIdQ26r+8tkRiY0ixkUK8I2le1Ac
Xf+GvLrMGEC80yn+l5IWn1o24r4If5XyvarpHrqdkcvjRgb9L5ZL/za16Bp5ayl/SkGL4GPiMDrY
BDdxC/1b5gzO6b1jqD0pe25l+MyvKOd5haJ8qG6ZE/8K1M8wCsCmePb8Crv7gG3OFkgPq0YWkrlr
cCeOmtYZiYZUb+xzCy7UWyfzwrFHz0UjWhK4sWpP8i3epMTEy4lec6MzWQVkU7cZecXM5vAFOJdB
WowUOGtYPnNv74Tx2CJ7eyAtlsO8vzMjvBuAjaSB7mcg9u5/YKW/ck/MbqH8OzngdE9NZpLzX92n
XHQlzoDOxudfqYMxhqOxJVSyhxrbt4PmesFw/9IbdUmsCx4X+V4AMIpB0tkhSjVil1u45524GhRV
wYfNPfZzGk/0cC6lO7Iei75WX14AZQdTlvgx5yNmSuyIbHfH/Yr9hBR9LBGgld6Gq63q805rHjqa
p5C2auCslTB+lYDnc6PH3ghw+jgL+GXgmSiqadnHRcoWnDC5bp4wvfD3TErKVyzyiVAas47mT3u6
0dNwdxPSG8G0AAfAKmnwaK/GQcE8pzPbyCNbQiEp1bfmxFKV3u6JLTjZzswAo+2fyNCD7xOdzZqh
Om7a3VJtk4CAE6BEw1aQFc+bLiHJnzLdsvSk85dARl1BikJh96iPDcfmQla34EWq0/UaZw38sSB1
ejsnw64vl6OFddNrHauWBC38wRCOLWFFKbm5ypp2JkgVNvehBOtkEFzH1DDvIF4DGMMIll9hNftC
BzDr+Bfm5h3U2gma7NLiqsp1OdXkKt7O+67nd9XyW+l9hY9hxprft485FP1f/nSyCZHV1JRs6Y1M
is6/dxf7t8IzJkRc0Kyhw/g1EJUf1fdm/7lGOgBkCCBQ9ZXeLFmc7XJp08oLKHCA6GGYz5+n63qy
942o5yGrBzm75tjfjnpYSkd2Pxo/bLFVS5pZuQj7aEK4FXnplt78FSM632j9aSVDhVSNvCEHT7uq
808PEqJE+zYK8NHIsdXIKHnPfml0fBBR/2c75hQ7+GS92EmsOkBXNHxajXtic0/dOjl+BF+ic0iM
1iKH33J7h9JBy970C5EFeOZ0XAQd1LpNnqQP7FbnAInQS75ZTJ2s/z5hkFmkH5xU3SDmdO4iVEDY
kjSu2mWV30X3ZT9flRSM71ksED3NvlhaH9CnZxTTvNJMDOlBVDvxwYhiOacHMnI55U1h8t68fVk3
5r+qhjFqfGlJnJ7o4OJWIJluvOZ8FdEWFpJKhAJcW0Yub5LrvPJxbcux4ACescjlkvBBKj4HwLV8
vokrOUOT+WLPf4hGWQgkCiDNp/D8mK/xnXL4t16JSJP75hr5y3bJLdg+yg2bqwZ5ALrJEL183AXE
rMcETX0+MkpN0DvMpeutRckyuL4lIJ6Ondk1WZpR0Ia18r30VeWotXyeork+ITyhuyY/tpE7VrG5
Gfwzm/uFrsGAyKWbB4KV6S841BXZQtZaA9h3ZJOFtMQfWiGoDHBWIGy6Bm99Er+xNjpvsBGfhNNS
F3fLj4PuCiBkYiVxU+gOmbCQ3UgQNBOvpnXcdefGmqdc30+xMS88EGh9oSLJzEC4RAtIu0VwHCp8
BTY4/dxwQI5OuMcS1KrYICd1z98j5plpMLvB0mBB8SZ1tVv+YRUFu9x+c57kdvjAZU1DG2rlXsDE
zYOyU/+hYpmiTvyVHnsX5ydMsDuUj+7XPncPMe7gokJon7w1eZnUJL1mW1mItu3fbIpZR7yN8d5d
bVZiXbDmMF1rCsKAyAIXv4inS3HZOHGhhfYVr+lYA2cs98CpnSiNg6VBR3Cg/eAX8Gc7q7JrJTLr
RsKkHQNwCg2mfK7ocTiywVB9KeklPv9gW8WxFsFp5ZSe5shyVNtKRGRVcJlDmLXGRP2RLGhf15nR
NqUbjtwMCjl02CMUroW9tIIf2IHZmjGiRVOgB/vWshhPFrGrGsOo8dS1OrTMV7wdx9cVXQ6gcKKX
3cK+UJiF8RoATEZgxMLYOGbjrdRD4LMRP9SJ5djaDHJuO23x0aGT5Xiz2rOfcvzUUBo396WbrrTG
G9meW9aiuq1Mp+wO/R9NzTyBdz8sCFaPuDceInYNWg6OwALJg/XOOK4pxNVYv9rzInk3XQcu1sqW
O6vvAL3zpKMdaYbRtRMJU+ZcQPBaoAWv0+T+Z/U0O1obNZxiE1KPOIgmQYFteKQcdAMZS3TUZ5Ac
1cG6n/1DPyCmHwa9se/B3hh+T6XZ5rfutH+Rcjg9GYskH0X8D430MUbev1j3jJV4ddEgIhnckour
ZduNWNaDrEHCgvVt5Fy8+MIVf4TS9J7p40Jv99HhHzusCStrdBkxVz8AlsZwqNlPX9XmHhiOBKTb
OfHVWVpVGSQ1VWUI83tgVBpqe390JZ8XAZWHIsI/vPYlFNUMx4MA3N336/3C9+IAXoQOcBnSt3KR
gLIHPY+TYAZPhaUmxjVQX1N1mQ/gU/ZveTPFSe/nK8C3QAxCE6KH8IJhuY5tM+awrLsZO0V5+Cc+
b+Ug0J5i40PFj848K70K+KgqAPq/tgkjK/c19zpug3GLHZDix+cKIOS7/vENsG04InKFTLnlxsbu
HlVTD3GxiY8hdvfNl4vQuFDg7+h9i7vGTNUAys9r3en7AMWyi3z30ywyud4PVxiXptf65LLGx9u4
3n2j7t9mhBhL26WQGvGl8ZB7uS561o7kIlHHNM2TiA8OBGagldmGdrXYgTohJ8EJexCy28gFAWWa
w5CojoEWOv70ZAS5axdWvAo4aGgmHnJPX+d3wo1SNWW9AABN5HnZNE7SppPSeNCLoiM+EARA7NdY
wdtUICZOciQ/UyOTlQQcNEm4Nq7Zrxq/vJsFE7tBRs2OaXTiyZjxDGkZIXVc7LgFB0Ao0sEJXqmK
KeMq4/wM9TtZpRKN4dKNfDga03aCAVh1NBM8URE7pmZmRx/1OVG0q0O2/Ko8O0RdSnkWDKzt2LCc
n9RedfKr3k+nZFECR7v1vzDoyaejSvo6BLt90PP5n2insxihLvpZr8dWLBJ4khCDovEghdvJ03e1
IOEpTi3ODjYWUQ3C3FRji8rhhDoY8Uc2rfdQmOJ5g+x0L4NP3lpApcPpuUh6ncyCnHVMeyYEFRWY
JT6ehXXXe+9Ff83dbtIN3xPeI5H0pU1aEUVa/LHdi7vW4IjQCVIGLKPCvgjwcwwKrJuS8pdeZIJF
fiZvMH4DI330M9QHa7Rso+ToYPxokCsQVqikx91T+eTamNozrhsiJDKTHrM3HOnOKeJ9WDvTTJzo
s4Et5M0o/VqjI34XYDp8M1P7fo+8P994VcvOOw21AhST4mVr6ekhtO/uLPc9qTP6uKq4HVLbLAAt
M1h/ZYIVt3Z7wtLO6WtF7twNPreSV19cxbDXl1I0wkrsHLPHeHxBLjy1vwWgulGWbUUHoM+DAOjo
TGrfZjNVUCu9ZooQ+LBtjUmbZIxfK/g/UOpoNS6LKpiSfinGGqMeSF/ltEudwGm8Qd2kwE8wIOOP
g5B4s1NLdoXqy2I/h2Cz68oukOpl4V9hziw0ntT0KDuKsfnuMHo8Rw2E6zKl2CRPyl4FDoZ9/h59
K/HBoR+Sy/Z/NDlscPyROSHWtIPkT+ta3gyu+tinTH4FPIlbRjeGSGjCcqorUQIbHs09CrqEOpr5
O2Jx5OZvxUg2zav1gOo48QQM6jl7NVRjd3h6hawyAy3MXdTS7q8QwTR3PB6DKkell2a0Yd5qBmBc
fr0ZeucfmzBFcL8kmxT6I4JHKxR3m2vS0hCst/v3d6IIxe2DxleQ95gFUJm/RYrDpYWLWuOT/cT2
53EXb6u6r+/HKD/hHmr0eopaLoLnm7g7rW6Ut99mwVVfZvo8DspS81pD0LlaSdzx4IiUA1R9Kf/8
em4j7NshzRfNLOmNYt5/wCSmtWr32URlfy2oaaU0bjyvLVMkJupqn+SVTimi2ixiVhWZZ6mtiZwI
SVadTh+Snax/ii74yI7btbrs9f41WdC5HZM5MBHTClblI2fn7EVfYJQKCmYK/rw9AB+smB6lUchh
q+SZO/HoTcBES3tBt2k7F7Phf5w9tcTONIy9VI5108/NLLG8bmuaUuuSDdPtiTaHAQmGw4spO7p2
CqSYgtLCC0MZ+1YP4RTXxRjefwE6Ohn396lKQj1r3ANmfF4sMdCZxgymZyHqwfXtcjx2vxVRiSNG
r7RZeR28BquChHFaU5jqKgUkOfaPCmuM/nwMQsT5PmjiTUk0yYbxHfgvXO4sKLZS4tPzls1y1HXl
O91uSbFB+ecKmwRvw2AKsfFgvxiFplb+GaUZhxSCNktIueCNweLzz3or6f0ipWHrnfo7EQl3Sqgg
5QTiTdIF5i0PZ0yKtpGNtbcb3rF3INiAeHPAP0j0z7Fyd8NxA9B2MEngEnucF3gEKVSMeasJDJek
E4y5E/ouM/RHL4Qcs6IanK984N/Ti6T6KEUqyMDFj7a/IH9YtRmvM8wpRYWV5XgZfZ0psTV9I+XT
03TriktRDjmECFq6Kf8K/ECGCxkMQ+kArLADkkSf+bE8b+WhWU9jDexl8KBhPW66VvmuogQS/jIm
1yhHUvp059sVf0DuMiuEN9x5vzC7C0FC4hAcZn0oc8uYnrvHNGRY7dofKNiTmYOYlvNSGAgI2iK3
cPtGupVetl/PTM3g7sEEGYWyMHK0V72NarkNSb4zqjIRZlBW+7uBrGItsToteufoI3+ehDE48YXb
GzCZSS4+mYLnnF/esBSC0Wl7te7EII5KlgMdkHbK1uShNS9vwt7aLYCFKBbti36A1DL2edahF84z
hC9oqWfvNi31AeZgSHn9iprqtoijNqOk0gmyFeptbNOX75BDxvHC7my8Bk6HVebxMEevQhIem1Ps
fbo46wnMEH1IdvJ6JV9AczUXC8R48yOZ0elWBSwaRpzSPyZucvpZ9e3Jrr3/PMRza5SBF8qStiGk
PJmxTvYk7fdPBCVCwtA/fEZtTAc5gkQiZ5X+StPK5P3sLQeVYBZp8GoSdMmq9Mv44/CJGNVW32xu
b+730IqXzE2bSniFamV215aqiydKujkpKx4rC1nSR9zL2sbo7W+uKllCRWdAlp6dx0RX9uglWZqI
DtZU9AbspUIpWJNISXrxZ7bK6N+Kqo07v7DYuWSWfkq5urpP4aNfAZs/D2ARMflKkd4Jz+n7lIBC
5zIpu4WCNlBCcD2NqxnTywINPRhxladTMTbxjhDMdERYugCt/4DKYww9Q1joL3IKcCyKjh4YM2Da
jrRs8Sp6NRqBjPnd6QQkgdLMbuAElChbJiDm/tTap2grG8GXruWf18z9PmtonBs/EvWRnYIkHMlf
yfKSV7DiIgQeJk20mwINRbExHlN5vLyXsI56AoLg0/q9E+l6mR1IvPj+u5lLsFMfGIaCqolNsj4k
UE2DDCOwXvToau7c7pFbD1icvw6ZJBPCpZ3aHNN1prMiEePKM2uH1gvBfFFWlDY+qD2+1mgpmceK
2bEMrT7itLuSBW3xJJgO+FIPqCtAWtuDaN7xSvoG1bIyg8eHMPb6HAo6r5GsNRFueE1KMs4M7tst
D4imsEj3eIibYVbEw/ESE5vbPM5XpH7nwssSGt0OLfBaDIZRnvYY5lY2SMlk3A+vIKaj6BfieTNb
CpZAonHQbbpaJJRkk1e+PDItjdgNDzP3eBBQzJgoQB8ChUgvqbf3UhfzE7h3fINIC3RPydWs0fd2
qaGu0g17SDFpvyi07TCI8/bYglxsPAm3p2XfSzCMe5PiUgHCxvJVUh0Uu9VmMjJ/YsmzQTmkkXdE
Fc+kZEsGjjmtn/Wze/LxvJgeA45ALQJatjHdNNlGLVM8YdlXoAJfLPq8pFoa0xuY268M/a2NJphH
6Z/N56L3jT1wnJY/1SBXITbUBi7L0zmsOBKNaT8VIHSub7Do1ziDOMUZWPksn1QiCvYEYnjVRmTA
1BVNd6BFmbFUHgJhj6pmiX3e5kobYIcGY9fwtWfQ/HshDRzlunfMnpaqDzpLC/K2V3+fdIX5vPGx
8DXoXccCARTgaVVhxIOVNAspM/nAvYNsy8d9YuOfOK6IbQ3iFbHCHZSIxttauv6818C4rtokNuBe
cTGNvkFo58AgR5hQk9B+hS/XxeVRZS4dcvbUY6Y8Dtpe269SrmrIDe71Wm5lUO0GP/5yNhsXpG+/
OOGmbsK5ljJSEwMjVj0EGEZStw5kw06DP9/e6t48h2T7wBC5PRA+j8Uxoozag8PeZ+HxUDC/hlBB
a5kZQTrUVAsU7I7Am7RrzZasPChgJZHFH0EuDUUca/tR7JcY8DH4/4/N33/3vHBav6NhrhHafWim
AwIf0Oo13XzoEhVpEywz4dxc7D+J7MoaRRXa4CB7zVg05789/9BM4IG5ruLTKgDZK+BpTV2Cb7PK
wCJ4kl/2T8imKirvcJcIWf5q4CRXHqkGse58sURLJiONlYLqRMsjL88S3aRYiYSQPbbWTiOto/oN
oKdPuoWJIskMHbC+ghg1l+vjdLWMY/amx07PGUCjSKL0CevsePHsAPp+OLw7wYOZRKawXw/UxuJr
4/WEyOStZdLUqxYFBfAx1BXiXyJUvmWITcn9VynDXbvSRRLwigta1vegkBB4/Qv5jLTsoeB7H1rR
8shDUq1zZaVchKQaRVj2EgF5vUyKy8FT2z8Fc6jbH26pAnV2mmKi8vnyu7u+8N5qlMqO7nBYncqE
mfDk3AYx/66OLal6yLfFbeYQ/VCj8teqQGxQ7bf1bQGQ2kIAgXfzXIqiNkYai26KuYSYK76OfI1O
3PjxUrFIyhhglIrbHgNe53tvz5d+W6Z/uG3hoHVHiyp13otYmjI4gsWmk9BJi4cSjPcxDVJ9jYZq
mlxiNZwU3sLh845seiAC/iUjOLGqhoSRnkzYw9cxJ4BtQb4xe6AiAWTMkWmUKNLQ+zazbitxBt3f
R26aeufG3uEd7aVKLJm49ZPz2eZotC3yirzBdOxtDMmkN2bzTlNJlNUpNwq759p+xnlFN8uV1o8k
1gdefZdm1chD6brIydOQOkGXDNeF0N/da1okUz8pgrRW7zavk1e0cJWPS4FV9wvqyGMppOD+x4AG
lP6KlYStg58BM/XKHmIe6GqQ3Wl0zDsJ1ikazwaygaoR7OtN/+jAyzly1t3CKg7dJy9+gaKmaBZS
x3MZqvQZ0zDtkBp7edx8m7J3rfZ0mcGNXwfpO0WJJUga1YGjkjCYLfphgmiCvABnpt61+bSq3okW
yXVSHBDMZO0Bf5suqiAsHTv0uijn3mGLQQURMXxlQHpSZ1duUZpPzY1lkzeRUBhsx7UFg/zNMZv0
LWHO3qLU1VEYk/+LcqGmKDxuDZUcFzJsCbWMA3eXJSsU7Uo/JWCr/5I3/FHBHLYQ7ZtySQInQjmJ
MW4D0PwIH/yjzbSKMh1c3YegrI094DcXAVs5TnXjSxlBLDCxjg7AymzokOwH4zZX9TyxypInSXxn
VJet2PrmhgaNqNKjtbv3Oztqxq1Aia91dQLOCjT9pDRYjdPoA+siJZyCWNofyTt3qJeNAa0qvEqO
AUOfEiezBnjz1g27ky67qzE8Orx7ACvi1zDS1JyCnEoEoQwa5X+oDfzJFH8ywAGz3bM+lr9HdW3R
wBGkMFJLd61X8t4qjVSamBMxli5I6yggnt20yyv5AO2uEIufOgDNqWs5JdVIIy4mcrbOcQ69F7nE
nlAiSYdvsscfS0U1EF58Q4dcXAjedtRJgFFKD0ONTAwnAfvLg1qc2FRTJL7fVVwgPInpOPXHW0iu
Fb3nGiJsKJ8fp07qwvmWU6GUGvR1GqwvtUimB4bUIyfi9s9SX29nc8ya2uRQcnM/NCW8ju9A8Dk5
WwOqA6PtHP8n5gzRIhrgrlnGukQsLhFKD9AdkZ8BERfhf2t3vLcEFOxZO/Mi5aLRdlcxJDOVLYi9
YrlsZCJPLFMe0XtMNT9jH9ds2MS+a2zOjIGeFi2QGrLhJI1rffZAFv7oVVTXRlvKTyInOMbzXDe3
xlgpDvwnaw1AdI09e7fzKslyRBQeW7e2yG3YOY20I6jQj5OTzNafVawsJYCF01f26fH4Zo/+KZfO
x/o/eOMxUQ+7rbp4+uZDus9HiKEvW3FMv/M8uB2OvzWDy0kjY6GZE7pMI54XPUbSOkqb5XSG2a1u
vNnQSbfkdv53RLXiDx9PJPAJgJnaxl8TOX6ZYXSRiXMcf+RE1g6p0J0sqxJT4xUU/n70j86EWuN/
+aWxZkySyLW+sE+lR2Ryo5toO+HxSc8XrCJms1zYLPvhsZhPP5cGyzrCaHHn2+3PzaAfIz+fWjz/
zl+D9v8MDtuEuF4k/SAyNPlFqhj8Rvcr+v3CdDMLSk4e7Y6DfYVgKcFjbdIjEfbkRAle6JmNX3EL
niaKd9y1II85hL0ZWiHhyfY4h7xKhekozeXV3P04laJCbOg16gD5IKCrPPgw9xEK5Yyzq7XbzQE7
QmfJg6mloVQqiRb85NxZC9IQDAv+Vp7sp3UG6uV1QZGafLpZR0DMvUGIQ/oz3UfJZZm4tbqKoOWZ
sm2NEerOsoty+vP0YlGXcJKD3rKXe2ek3Q62wSo1DDFp5cLXZo4xDDrXcKQmfrjq5djwlETOODDp
YN/WDC4BkOWfB4mhbNrwyHPJaknHAcBHygQtqYDypQ2eVtV1LbDDYqRKoGdHmOurWmL2ITBWW6Gv
FGXPjWqgJd6LNw+R1Jj2XIaH3te2unR+EFjlM5yawL9MzCW9k2ROmDNfpKAHx20ro82KEYixf9ki
MMfoKDw/kkzo1dX9z3KQV7imSFc9HLlzLRgPNr4q7o9U94JAI7Njdp9GHqQJ9rULwvTyLgZfSo/9
g4s+vlih8r2tfDj3Gyabl28zbHQcINSTIgSUAp/jEM6+3W89gIFbrp44yOje5MeXHwZOcBHx1IFX
skW7nxVZdd/LtrqU++q1zFMJh3cXePjCFIWoG+olPa5AD/A2TjzTxEti6ctj6Qa7JS/ILr0ixR0J
ZZLO/7hcp4xXjOzkH4n0I9YL1jXDZ6Q7hI/VvJwrNXYWVqeSPqJYkC9a9h7XeOJ1NIxrlcR49Xbb
EXv5RxPTwvhSi6sDteT4Prep2vPAgfgW05hGeXPHP1iDxbfjAOSTnwYJhOHAldXLGiHofxSUNX86
a0jntvaXent0i0mzd8+5m6vrLBzXXVO/P+FiLCYIUEY3hEpbDIfo/nmg0RYxL6O7EoMRFwh6ZDNR
0k79ojdpGWooU9OoZr3yI5TYE/nh8X2SIrA27qDEGat1VKlytzxKcLMNklPnpaoeuiIvA7ZddKaC
2Qpip/hg9A9XfLLcK0wESVxHrs95LuPxQvkaorNBockd5ybeKDvucdwCM9F1+vntNO/0rHiEFbun
4xKWbuD2W4kDtVzXiWM7H5mJHmPLaE0akazKWfJ/LJ51cOmllWvxokDSdkzKgYi3P31EzWKvg1XK
etprtz3mayeIv7jhG2l0wvV/bx3HfIFDsuZjxwH1IE82ErWbKRFywByGif7nGlNvXOo8o16pjLec
9/vtcUXOvTUXdpU+UCvkQebJbTyfSmkdoG4sq1GgWgMOgg9mu69j3bxnX6tH6DuHMHsk+vdySf1l
pqoBBTqodXP0wXZepesgnxIKrfftT5DdYHb31RICk0bubZhv1285nPwmxC3Ho9iuhbaEsATOZ51i
EQ1gL+zpWD9OJSamQBFaCtClrFR33dwraUI/VIlwVUMm7ZhzMTQltKFwhnIMNCBBrPm0sPsGVBvk
MYTY6u0McIBjEtnvTrxBD6liIWCppKI4E2yzuPu6RUlST0Wif2t/QfV8BXg748w6YJoVLwaMq97N
EEaoz03C1/dquGVrDjfTLgEid7b86CuGnqozTT3fscXVNFt1+cncM119DNlbpcc+xOQkapMVrmFG
SaAzP8COIIPvivj6htjmj+ptYbp44lru970d8lPj9VGSxo8VPP7WT3rkwPN8f7OqK3X8ONfcPzJ5
+fOJmS5MNcGDLdR9ToXQEIQT+lMugCGZkL6Nl0QzgmzSpd2ESlskvi3W/pbAF80kCCo5REYt9f2b
8Ma+JjrkwTISLm0WbdewEigGJSD8f1fU/qLuLTMmap7TUz9KvxyrE5SV9iKs2XiecDhVO/TO38yl
9Bj0Wa6DwiaItI84Ghz3S1wP8X51aYmhd7tyUKsb/Labk3c2fCbLKkqH328zlt4DqLj4wl2iGDzg
qkgWMVB3HeB5vtKvPL3M/DipHq67cT4WE3VTb0DKXUgtHLpfEZzXdW9UUuGN7Tu4VDEjcNmjycUU
+vBWMErGk15Kq4dvf3NIRyRcqoDqm75o/UB1TUKLYe0ukrQ1dNnDoBSGsQaIr0LZCzQmwPTtqynJ
UzjRzjFDNT5p7p5CN6pgbiaqTEc6TUN2AzPSrNko3s6qSPL6ay0KpJmY0efQri1Si2veZqAZYEH4
W1BU5IAuSmClU84yMbRFHa5NG4guI+t5LOqDrhYxAgnF2Fz7iwV4Yz/qJcqiHAm7AFPc/p5zg7Ms
pLkVbnfiUoIZzAKsZ5+9qt3uTXQvpw3F/3n02zfPAXje2lVg+VccfSkxKWIF8pMtyEhbHfR3zRSu
RXqPoe7cQqC9u9fPW2LDEy0QliAon2owVJA24mD6u0F0kkURoXfQ9ww6ndD4WsKoDkxIqs/lSuCv
U/Wl5OCYGZSQgFc6V+qILY3gGs7iThNcujfvnR5if7MrWY768riWLzR0sNWRdKYs6nRpqbpvbvoH
N5SROUmpE3U81l4xfZpcUDTONN3o+jfGb+Wmy8FAqujxVYV007M+N1X6diU0TiZowWVaHWWR36NC
Zg58ozYXaS/o6r+XCxk7RyY78ZjJ0Xg57CTOgxFMggwVJXjyE1Xh3aCvKPe8L0BNl3YEvlAfNIlj
KVqDASxhAqaKS88KstFt9NElKUp7392a1hoYLYsetZ9kHKFX//3jdUpUjNZsp9X7obHtBe5H7IS+
Ut9hai9EK2bUVVF9eS94s6na4PHfd1wfpDlzGM0KQuaoDuBCSCDISP/Bmq/zm9XfpCZnMzKdgy8h
1f5Iq1wcsFwMQctiOse3uLT+zaHwo6uxbwGloDDqfUbatypy8zd11l6ukCodnEZ2j7sELSuGMd5g
Shpg9p0RTC2U5L1aOGjRVAq0IHKd7bMdD/yHU2MwoPeDQGWfm4EW0AEQCh76y0AhFlpOLE016WJg
Tx95Tr5zvWwOkV1ZQqw8omyXdaG0o5WufWepOCOGROYQ7DCY8TzeA3mSyYNw8WQ8C7Q1MqaCfWbT
4nmEABsBxjB2xTGp4q4s9wP89R1yg3Xti11h+msrdZLoqDyVlyR6r+7E1dZYqWccZdWiATmjHaoW
H5iP8Aoai1jRs89NKBQbDxJoIZycHLiWdKezCUWw9TCvfek0OHKtmJ5weMgSwvqiWKmkqKTmJto2
4LK50xMH4Df07oLhLqlnAtOs8ansO3SDoJMb70T9Yn70VtnfuEGzG9Pz2MbZkVs41TzY1K6TBpCq
oOc/HlgFttNMQNts3qAbzcSXHfI9giDp7TeTm/uCeHcxYJrcevR/QyAVEzBRTch4r3x+z5lz9eH1
eOM2rd0iMBSpW+AhjYc3T41tn2HEpzlUKNOJRJMP+bDDOaL2Iw5ftl0lqq2K6OIEgGvGNEkRLqar
eGiXvXO2rOV54dRCEEIKBRudDJ+MuQ3xC/FCxG7JHpmYHgUQhziqO9lE9ZkN7V/otjHkmIIhCCdL
/fHV6BMWvxTwV9zMA8bqvtEK0/h+LL7ckoLZqgV9pxyaIB3bnJ7EtbqICHE+F0/XAtIIqgfSJ6QV
Ghao6XdQA00gnjRwYNO7VbY+rohPYPOfPExPO9TXusbCCPPF00XDi5KjtxUzq1VJendlbKrdIHaO
C5/QvCagTEqb/qOEJBvjBYEh4j8Zq6RtUnpiBPJ0abYGG7gOy/NHNY0qzaOa9zsSmYXPAKjawYPj
YHH5XqAnHpLM46HG2lScMJsKBDPOPoXh4wsQdfS+TV3NhdotHgF87kuFtO2iaFCRldZFYSqDRtmH
wDyBlwAZEqjdAh9sSifXNx9GYgO+Ohcjn25hAbNDNVHvyFJxOT/0cYY7d1YXAVYi5YrRZEVF+R72
oxpQPmlEwabxK/K7MIglcpU2YgVvGraVZ3f1cfHscamadN2Az6afVRjSHZYsncxlsiPfk+5GUB3p
ouvAiQA+jEDJUrYrfEqJ3HYw1zshGLt7nstGfd9aFXQf+fWVSeeGXK1E5vJ1n7EPK18YSRt4diN6
+rS495V9DEyF1e1wJlcjmQZlIfa2BDH1fMXBGLqUPFV7o2nUF7HZYuGO8b+MaawemOYOD+ZS10vt
cI4TaklUyMoabPXHv05RDeAB7XTDYXNgAfVf6EDI2nW3MDMWkr0uXTiGzGVfXxvoZAQBFZPpIdb5
NEWiwduMe8RLXo3W+Zv8V88NXx3f4g7cc5gIzzFT/sEiw/iP+MX9V7dYj7LYi6Tl5n+4tFv0Zjhg
AnntRKT2ss1YXFwdpZdvcZgvHV9kvALmNLkcZDQMJYe2MkPwgUX2yXlXdUOO+YiqhBmZx8PiaO26
PXHuT3QZ6NoThc1uqq12FrsJccG3EPlT7+jEnXDMPBKsw0MjJisk6oLTxPeObCQ/SPhcOZxe4kg3
u3odHgW9kgDz5KCuUFUTRj8yHO0VNtvjwB0yWVuycJPtpOjNMQIJ8HSP0H7Kk9zruuP0I+KVle4E
zHUvpJj4P0+QcTIXU625wt9OOtuMZmLBqpzNoUeLorshtuLp2qcIaiOOGaULeP2RfoiJnZU5QChN
ar1U/foWcKsfC7lwX24bMv6ZII4nLob6/YTktid5h9aOLXUKGFKaad2dX5Yz3mC1yJu4yScEx5Bk
iZ5WUmHP39GkuMzWqm9V3GUf00UDC3EDSMaS3UEJVu2EwCNIYOv+grVdFZ29S4muwrPBi55kU/lS
mkC88R25Px5Rgs8Wz90TDVHgdHFv4PCvfQ2jhbxUS4QtjpBRPkj1GmoxS6k67ukggh3RudEuBCMh
f0D7QaXWqbHz49nvSVB34zh4681Lr73SQF59dcrt/dyanvDGpIJbm0oVfZ/ZROsmDRFfmoLII70O
zqu/xmVZrCdXAjOK30A49pZVvpvYosvaTO4cxoOd1fU3OB74JR83jHydfr5DIwxSKCN706FLSMfK
wCOoDdiwNPDabtQddA6waTTry5P9CbcyKp+Ia5ngmnJyWljsW16VUFc/PRV8t6ARyAC2KgZ0qF/t
Kd1bldfkLAM02UGISvTVA8e9Q6KMnhc8sD6YHVE1eAmrs09eyN81JTW4fGLPgmhBme3WAsSDTs7U
tJtTutjLjy3tMDmtpTxsq2HYG2c9If2Xg7VZFZ3fEHU2GzX95IdTZ6nayPVP6rpLTWHAN7sz6LiL
zatKVInStH5+4F/1uRZWRDL688+TexhnWrimG/AJLCWmKE5u02vMKDj+nrNj53ee2/bkBuc2BX+K
b77By137KC6ThTojdRaNltRh+Kw+XYnm9yV6X+w45tb9J1f6/heVowpFuWPmtLeq1OSLEpFbBZyW
c4lYd3gJVh8nwbFRcYYiEXqgDzz8rZMAQKY09/NccId7Ij6qdPOJ75P9HznFcLOR9k+TSOEK2bMa
uAwMDbrhCVsmXD1jI2DMne1r7Jp6kL34xzRQLuhLfvUydYKFeFpIGSJQEyFUFhftX2N1JpwNO82u
1X9DTDjuJ7fd4rOnJB6FbjZivbvp8sjwxzmuSjdT5qBnE9z8WthQ5jB4dtp3Xw/sXTs1qxlmUwOX
k+ddgndZl5ngGzxfXFlj3A3xIqCrDgTuYzarA+I+zGvG3wjprK3i8nC6uwC9IDF4Ddo6OxhRBRfl
bmA8flDyUdYs4w4f6SoEhWvh7OuUaAD906b2Y1gQGGjRjtA1ma+i3LP75a79fYcZW8FgSBayRRdf
CmRu4eiWRqq8k5rpSDZsFjE6G5P5iGyQPn/68Eq3J6Axf5EbUSE78VWF7bTlEplS3zThgKHKnGEs
GdqPye2arQdmwcwRWBIlyz4cggmJk47eVo8QIQ0CDu4XQ15+fALpl+hA6GWdFAF7HaCZR7+P1tD+
LN6PWe2HPkmHXgafjNtItTVPf0j49hcxd2UWrwL6wgA6g4n1aX7btBYVpwH92aVkk9uPw3iabKyN
mWOwEVJpI+mfNZN26MbqyK1KsUPBUa78FIYGTDqocsayyYXVgdtK5R0hv71Lh2kgO70bnuzYkDzU
0NzIysop09z/5v/2gZdRnibVTKM2tyCJbr0UE6J0hUeGFCl0yRFaowXIZ+eWxfEyfimEMJ979k7D
AEdlTowndmdd+IMm5nZnWa1A9E+6oFNEBujv95Ia4kfCyCUfUCW4tz2Qictdf7MZW+hqD61G51G/
2IDzv0Lj16dbqsgNQAGIF4T+QrsOlFCgd9qT7iJCTLgvktd00osutaS2iYEINxg2FARlWEWyBSc1
8hY8mWsTYFQpH94/8a9AIkJXinomUtWC7faBXOocp0FjWlmxDjmMmH7rQj4+68QIOU6CItCS2m7c
SANsqe9YRzPSQmLViLofv9CFJd2/zph9fz339uOpVIJtCHyR1ybXneiXSb6B6JnX7Bd3YmBcyJ36
cW1DLoFIu1n1PTrHZyZYdr+rjnC5pZIrli2m9zXlm2J4v5nwv5/FHeUxbOGauKElWC5gtgssOtZG
XDKgRojGL28xsISQYwhAHrIkgnG39/6Iv54MgmJEtE4fII+xcpNozKgGW3d3QGA5LzKkJdfwn97U
6f+hc1+JH6EWzrVAsp68P1Rw/q/lh2fjNdltwaVCfoYs6AgjBq5/ZIgCWhMwb0vh20Z8CVlhhNTE
blsDl06tSgQ357WhRfMvVMThzW8WQ8mLvChDvlmo1aD4ysmy2hZZJRY347AO2AlFjh65OckEVsKa
XbEFiSZdKx3bvpFcYSg4MFs7V3gXUkyR4eTOcLGEXSemhSIeEpA9v6NsUTzylVse4+7onXVWOTpr
X6GgWUPk+xtHhTzKisqYZl8s0EkpdAvTnX5XgClXmHoPrXHeA6AnI+tP3tlgSJZ2yjD2hcA1GNG9
eosfwwwAJ1xPcUpwlW/Xtf1doyw9ph9vkAOGcDEHnvV4sCFgvS0xNVwvlGj6auL6MbptIqLeqodZ
OanDOOI6lxrqG1bfmAjVZf/+iXy4biB5sWRBbmOzeXG28tKRpZzOb6zIfL8NaCYxuGHoVTVZQtah
bNLq9OlJoZHjQLA1xaAopdCbkV56YTaGspikLrYAHGyMoy+i/jOjxs6f9RO+z8C8BsM82npda9Vd
GUZpb8B+wdadHDqh85v5kLzi3leXoXjlYXZzmYykjyZuKno83Irp31taOhwpw0UrH9jANwZ3GihH
egg1ra2Eaid+CWa9vBBASnsQb2TjF6eeg9HlR0vzHjrRKKGF96V1qMgrYbeppRH974QcHutcFBsi
8gnirOSvBQ20k50oFqHNXpaQlTopt1s1Y4zGPEytWQYHfIQ79DRT8DKdWshBWKm8QrxkTdGgNBZb
1drE1wUqYUFBolheqHr0hDBsxitVyvUOh/pw3JdodTrFrrnfTNB/7R54PTmeyX3RfcmXyW072unN
1QrW8uNvmplqSUWkHL+3FJobmG9pxda2uHYb+uU0PfYSVGhEdtfwax7zylESnO4ZHtDC1PorRCdx
j6dhdFrOthIfYf3/N+8wfEKYUSNwi3Gu8dA7l6qSEbRLgx9iUeYDbNKyXLwEddQpVwa13RCQPGGD
XcZy1sOvYanud3kicvJqViuH/QnqQ2gwIA5huH9NlBM7oGml4Bu0G7i/IU25P7WUSOtSBk4Mvwaa
r6t2pPcH1/qW2wH1W3yACyeeu3xDoQLlv3hL7AwXRnF0DWov6lq8CnX8R4BegFkuOpZonLSc+k8y
EeIAkj9ZRGnATbM5JIW5qQW7NWDkCM/Whlx0xYgqIh27rgi74iV5meYBwIvN8tQ+LUmFjJHb955k
NE+O61Bek5Y3GHr+kxaj4zUjq1OgHak1X8mDfkvhVJIabiyfexYrJxzORNN6pTcuu5KOF+RDE0SA
n4/mVOgXmiVVzUrogpPdb46gRHwo88TP9It/U3rKmEK/PcME2EngxtnwZDt3lcCHixz6bdXI51Og
eVjwJIXjHQPl9sxWTzHvBBPVOy66RW5lecOZLGw3umJNpu1UXA5xFsy3+BI1Dr7ZH/Q79M7cWsjO
ADf/k322YqT0LP6rzhN6V9GlwHznnkuE3hQjzGvCbTHIiLBCMmtjCsvth+zE0lKBukBlmKBky+Ac
smzDFSXiX+YgQLMFxhCwp1qTGz0XnnrzH9UtTszQaqDLMYD/sGVzxetryQStKd0e/Zcz14uQJzi5
RyQSMPXnLOuWsTYGuer6BgKvEmBMVy2FsDyg4XDdB6B7u0HjPF5bfQ3FfxRiX/E8gxFyUm6nocN4
wWq+fedNIZMOq2pDd4r1lL9FntBux/Q1bfSC5roBLFKMxucASiDxFlCcp3EyDDj2oUgAUTeOgbiO
FnL655SsDJJEqcZZWLbDad7oI3RGCETx2GmI1NfIdVUV5bPIcnxve0et+m1No4Hm/nyiB4vYMAJI
OWhf9DSb2sKm7+LQDAlz6fua2Q5EvKgtyxCTL7RDgtqtg1OMrcpMFOPxroo8/0NNx+lub1jjfcBl
vCB1XkwgNvSfT0YWCHbwdMW/f+z0HoIgmkFmAVvQNsa3dY4JmoiiSHIq1GRmIlyIgxbRRdOQeaQ8
lyPU7drco2WEqKaNzNjoePmPolIu/3rtqHhtpOdbAqRiOLEn8jxDLGpEUc7ODgKLaKqzWY+8aYtb
cmLqs0ogNMFyj6+KB7OJINiHx/8/L2qXVS/pRaM625J/LWhtSO+0Co5QtvzYe+3PV6hKrD1tQPEc
Xs2N+Ka6HDAyO6FfzOWvAS8KsmTnYuCDHfgFgxMNAgwdv/rIFkHZfoxK7cIapQjcllwjKRv/MZXE
Y+3TfyJ91vrivld0y/ysu3THK97mnpNZnF1T9b1Ey7CgJvhQdCjHjNb2B9p8RMRspfFv30OgQkyP
JurUvCosuGcYVAXDGXpK0UW23e1HCW5aZNRYepRSAXdXtHu6666zlmNavqWLHT8bEh+bVpWczn5T
gDkYj+Vme1ptRvy1JinB3S6mjvW37VzkGukS3ulXQvdzZXyHi9YTozr1Z6QL+71LHsjar1VGuF1f
hBx8veo89sQjBDqD++o17y+Z3WAOIqmlKG0f23rkGb/5nGoGQJmmcwW3dGxMPlb9pRlCzeg+lvwa
tmBEQEvulksQWOYt7goo5xbQDUmu7F7v2DQGEGJooEj/LWJ2KVqdW2ngPbwvm39uDRZHdeWB19TA
tHCWN58Fga25uYES3We82VJhlM/vmVVjw8rg1bjEESX9TwR2zgFsuHgH+Vy3ScwxPY22leveojln
FeLyf+vw3jQAUd//w/PHeF9Ua822j/zid8e4R+JCbEr/DJuAw4/1uuhf4LcI6AyP2PYZ/fmBpaFw
0ZzbwqQ/7vQRR+/h9zDFYPTV8TFQIZsNaKB4AvBZK/oMDLdD4d1LVaiNHDZByVR0YLE/Ol3TZ8LJ
ZqqWyUi876JLY8zTV0n2DVoUihYnyrprwijzFlVdym8d5uOZdnLJ7ANehjT1+jf2bTbG9uzL+gL3
mMWxSJbWDl9I4/rtg5gyoHysCjLNxV6x6lvg8nMKSpxqemhsIz5y8ZpE7KOd8jerJtUmzXyuvAZY
1NpoGcKN0VKdCAoo2kYDczpNlJTSHMk0/mg0XmqxbAEI5/yKRKD282u/cIdmExX10bGRBgzg7lwo
awjyQimUHqu33hNZVXt3NMduR22K0WVzqWj79RLKrCBSMu5EpeFtgOqyshuyo+pGKIwoDhR6bg8T
pUv+L3Djbx4XRiQka5g08locvDbQaJtBEthImNXDD3gvNcRIwRcrjxZrY/55JMrqPKqfCHVkYGAy
OlcgOuziJs2/DBdnhox2JziV331tSaUMvHE+obC90evfbj5YpSUik6JHwfrC8Uc9Pk74M8xAItSz
qNkeRitoqjn3YhN7ldXgzCWUF5nQw+uwhsikuiNZVHsBMYY+OCT7mDgTDt21cIpyyEvVowpp19Im
/B4UB8bgfJ6aTDJT2eBh6RbTE48tjqWnJIChCwX2IgISElPykiH6cFgAHWGN+9u2TlWmy45+nrjN
em2yVpcO+LowCNY46qfxe41sl676l3xqQsJr3tkwHOUX3NTRy24tznPfzew+xORfjAik9WQt4vfD
kK5msMxWzGzrBzKY3c5LQ3ecWNsuw7WrNJmiWvUbephV7lc0U9ML2n5tTwoSdvxRBFK1G4yCFRnV
ey/wUjq6IHW20qH9QujnQo4HhdEf35BCP/bdsMOOHItHGHQwG+6D/QvNVKAK3J+fvx0OyLd89Xxt
6KHmCLiCw4Ra44VMU+TySPZrhCWrfeIhR4Iy1FFz4BdziOqxQhzU+erDQFAjH5jyracZnzAF4gfD
AERlpGhrEIhxvZLHhc5E9XBB1f4PxiwLIDuJWN1b2ewNbEzYorbDhLHH3uskSBFLWUQJKvJv0s72
j0iYVx3ndlSfg5ENispseH99MhE+yaeMoHPm+wRU1VrnD+X4eaDDctPSX+odK5ZdHJRrD0St6Lie
bQlu7RaC71jc45mz7QpkySsOOENPGUJIh52mY9ddD0PRRNNNm/w+Z3f9bi5Y0i66PrhgULbnkW7W
PU+cGtULNSJGfwZ2Eac4tqxPfdRXJ7JxSQ9EQ9oJcA+RQinYoJ914H472fwMpoRwjPGmk5nrJwTI
hbNX+ucknYI3fAqtFwMIaRsZOXfUws6D8T7Ux6R0W5LTH6f8LzQOyE73psNdWHETYv7oYrCNfUM/
7FvYovhGepl6t9oS7tOEIfKWNb38PjR/Y684XkDt1VyGTs4rokyCBX/Ab34BXEUa/xe+L7FpSe9U
Ew09Z37ODqP4NeWYQhAOBzG3Ee8AWf/cctb/fdaiB3Wi3xEOH16KC/FGZ3HvSpoZrqU9VNsr5MIc
mYdEm9vD9Wj2CB7VKxFpf0fJ+9WgHzbMXg/KluGoEpWKvVVLCuALGnK8WVhKQmmof+tnzHp4K+jj
tmQmk7jQ/+B7f+wMg9QgN1nqAMS41LP1B1WuS2fydOSWiMiAJM9Cx9hC3qGeV12AhA3JGiMw0Ew2
PpSBCprZ9qftwRYsPxoDvNC7bNFiD5xhwuMXS5uk4+7eWUWEiciubmnjhNCR2jX7I0a8eFoMF2EH
WNHFDAPU3Fr4C/ay09e/pDTH0x5ZFXdQl6g3o/TPk9+MXr/vH00l5njNneNIAiddG2GyA+KWJBDS
BHQoaZTZDIi7RqY0bvme2PEaRskoJqEJMJ9R8sZSmQtfdWE1gCymXzdIiCby2zMNcUko3g/+cFGw
78TmJoBMbJnIxNqc+uAGHbhtU0dnHb8cCJMuti/67v1TyvlLGeL+UHsJ3UQNx/DFdHYRHpQ8Hl6o
rjCkju2IxcQAC+KJk9o6PMHM40O3kgSo5p1A9G8mSiimINbMJwdCYxNC0bHE8ryt3tiiH2uV1BSb
w6YV69WzpByRA2X6q50bG5nYVYoYKXvgENAc8HYdZptJz3wC/f/bp+Kmb0I9lS+DbwCDS1RiqezW
KO7KA4aWbddYd/ixt3mojVs7mYdllf+gsS6YZiSNhU86oBx4/C4Zd/uKTLEga8YkyIGIEQpZlvJq
Le1WyyQvEP2b50KDhDNObYZ5KPVfiE3ZoVMRO1Iv9l/ccL5WuSwWG/aJgg7DItwUNry9QvG8liX1
2Kj7Xpsu4P2e5PWCb7+zkKRa/aza30DeV/xgmV+3VaH8jomDB/D2ZSVHNnuwePIDUMGXV8nWG47w
3A1KSJNnCEM0joQtCVjRmQZr1rR9j8GQOz2RDj1sX/x4l5h3y87wIx4F/EajAG2A0aGiYX+JUsOs
sQXq8P/FcKFb6s66W36PN58uBu0WcszlvXa/YkJcbI7pz9YQdQh8mlQ31lLhOiYFGUxkoBoUfIK+
46oKh8DdxnUBZdD3Y3ndivIjj7tc1KpJ31HeCoIDlmnC6XFDl8C/gCRKWr24POQcBc0MWTr4GS9R
zsx4kLouqDhc+rBLWPvqo5wgb8ngOTtoOxKUhyVaWg55UAz29mvJpD+9Oe/CN98MQWZHdWqay2Fe
sJJNoYaoafcsHnlmx6byXXndKSHzaLdfHWXY+huoDORuOipOS0E5Grc45lcJDmzdsNpWc+fpD5QP
7L48bJSzcwVr51TCAtN6N3aByRLWMNbG5vjrJ7e6fz3fNkjVDo/YXlXY+nAyjaz8BexIx9Sat2l8
38rduhUY+/hVW/dOapb3xINdtFBY78gu14oVr9/mvU5yyp1dLHMvrcPW6VsJaODDnnimTlehwoSo
670oP6E4lHi3MW6dEKDqwJjD5MUTPWMqm8yZ2KmzjszCL6PA13kmpRETrPwJXodboyOzLgSUG+gU
fJWfRb6q7NTik5V1TCsc+kW4jEUHcmno1WDNbDRtiiLU+QJ2oIhT88Cmbh4GeDOCtVIFanNA+kOR
OwWX8sfD/vmRw7qCSHPEyYfqRI5S8TmmC5hKHNfeZZeLJ5Yf6WSR6MYH0/cEN6qs+smh+HhnrSBx
6vTgNrqCoMjZv6pr8YwcNLH4U09q0tjL84t0CcTZFtu42gbQas+xBzF8lSlmZL3aedUfDOlUqGno
xgrEc6uxm19S4kABv6Cc0IxscYGbBNJFPvO7w+gm22IlpfhwbBcxCQR5bH25Zjdpx6w48B0n7Iaa
6Yhu8mzZcCCidKjOFI8KHvQWT9UY7blHd2EG98aJhgTXc0kCRimOMRnQmNWWDayDui89LH/15V9y
EqMGzrMJ0Ok9xnDwhwdmqQdKIqA86HL6+Kf1jUmMl38kfTkFdFOovmyE7TKcsrx2IBaOd1za/yip
1/OfSSrlC8tjcEJaoiUs/zYjASUKCOFQtINeaX56F8SpHGgvwazzvupfaA2shXRCaVTW7w1KwwMz
g7CPa4blAciPI7zp81ENUnF1zHnQeymTEz1g/cAoRnnzpNVtqr0qBlOVgvw4K58PSb0eyFvLz9D5
mSCck5VPdW8KbW/fnvQJShme5WF67mVnuJCQq5aRmWHwlI5HUKbnzySC05zrMkdCg4ojEyt4RQGU
kVtjUys7dx/nr3bCBIA88AsMe4r84eAfPOrXaEQ38LfcvRLNQWGBVLMBYMFhQATyVLA7jnIOvNzy
SPEwH0VaCALIDy9UOdeo6mnHVUnH/W5Ud5uXM1zxt/sSS+ZHl4dwfEhPD3H5275ChbhGxC6HHbLV
ulsYEJLrT3uqXFKvpBNXUXufwf1D4BEq5hpvOO0lEB3sQZc8hjjX/RxefmZd34BMN4/XuppYNtBx
/oxGtRAYO3VfheyBZcada+z7G+jMR57AJYX/mszn0P3E9d5+GdZMqRjeR0jH9i4q5ydah0rsrg70
+Naxopk2uh+Gk8o5mhQ/NrE3ZRFiPdqZ+7vXfHucbbNSdXbdSggR/p+j8nDEWDeAo0ZN/F0ddm0C
mTOVkzpb+uqQDubvqfAHI8MdwMoHSDTOVA1HiTqatzhuW76hKIF9yDIVWvY95fwz9Xz07k7eX2N5
5FKE68P6JwgXUTWioZy8qXCMizqDTimQbdivQQ4wiiHGCL9xoMvTO0/XiEpE+KP68GbJf1p0DLxM
SgZdyxBbmYg8uPr8vnnXVOjvZD1gR8OTKEWbTFGxNLbrg874r2flvhou1NrWNOmoVFsUuryH7qGb
geICoyCCAsMbCNcoPHBqwkgJUAkr59KUakqH4f1Hd3nJaxrynVnh636fZ1swl57n2Y+1f8onccCH
qX3+v1WzonO+X2fKCTtBrV5kx96NZrgu7w//NLgVvWMXss7iC2eKEI/bNH9xe/xuGGuVn2hDke8z
23UU6CUe//tl8KoWL9gMZSGcg+YRB9JtS8bI+PLjy4btOTrcOS2POAt0rjuN7INK4cNWYBzJGTX2
lCI+UxxL59ptydeem+yLLosDJrmP8CsJdFYB/eF2ucsAAe/n7jT7E/4+imuCJoWmjWoLniYW0z2l
rrAq57FvwSwVaDHxvxZOuO7hOFEB5BaQ97viRzFEYVekrDzgcPbZmPWB9CnX/oPirT5pJN2aIt4l
h4Gr+ms+FnVsKfE5BC+PL+Azv4vFw1KrJ0TN0uxMvWtekb79bkflf5IGYmn6O/v/OAK0Q6WhKZqo
feqjPwzEBoSSbes1eI18Wf1UtTCbfZY/bZzzFYvYjPB/gFKEfDyl6cSUtkpFZyCSJHFqbrqFD2N/
rWtlnfbYLG8Mu4++zLgEtDhYGcWxPDOB1PoOSivi1s/OPAFXX/Nx2woYSMrt6pXOHz2+X4DwnDjP
J0qS7JIMg/+L5x3zzi+ZC4IbSpibUpeageJNM2G91OUsfWchrhsrjK8wFwFuZ7TRkTh1PlOp88K1
n2GlC8HD7fNL0md33//upKuMYqlQ4L5WNIhy2/meWzYKtTeFue5k6eGsIXoNcJW6owDiVsYL+kDD
IZIYWZaI8hOzKXjWQZEZVK27CNo7Zm+WKQHT/rF2pFA95bslegLyXjOdyQam19UckTTQMTaiBkT6
+8srVkw9uLnNgG6oxsqeeC1DgbACHj+L8KART+c/w2pl99JAtpdVTNuyMdhzzpvhkizwkQtA0Yz3
3St/2sdUmPMCr5Q2se2UBo4SkmqipkZXotu4F7juyLMTKLixiARqdczfQjptxoE3hZ9o0sEe+JFy
zpp55sjhgtnpx861nNpU7z1TxdJUZAZO79/aDD2aOM3wc9efRc6Oi66ZufdN+heOdJCuM/Ebi63b
aYWIBHLE/oIAGASwtOslQjnc+OVOcDZZmTmW9lkODgMn/KVo/kz20lqwQOqTgLVOoUBJP1b57zEO
jrm+l2WURtZjHjnrjTfAA9IM+m1ADEpoaoNXPB3CWtHCgP+dQBeTrim8JKcJgP2y9QPv6XkCiz0z
OlpsKfwIgH65GiUgnBOQ6I8W5HFeOv0vV9yYNWIrlcCHKgHmYNY3tV54kRf60Vgsoji7x8n1a6hb
pjtHi1mFHn2yfeX4+YsZKKEyUkEyygkygnfc3+TrFJGlh+D2/SvQUiC9L7bFlWIQP1ICWBi05Mr+
gNfVhAtEbKSGqFAz2ibYtKSNgcURMGBez7t5QGLP7f4MI40pSkABRmayDWqTGBM81QLS9u1YaBV1
g88bjcOQMVRaAcvCxfda/ywWAogURfJyTrlWWN4YJNIWvrI5YF9uL7ILiJ93h615OACtqrj5n9Vk
z/X0kh9gqw9ns4uvXzp3UPLRNG812QR/N9QAiq+3JLCpaNZJMJ43ipgWR0mb8Q4jCn22+6v6Cw7T
6vFoPUAEsG4DmgpuR/3io2CmwfZ6pZ3RHDr1V7/BoRUUYn/Q+XUNmlmHD5cDP9eJ2GAiZ3PKYAg/
jGTZiWmm3kSZ9/tsbCN/PJsI+RVYu5eY64nGCbyywKBRaAkycx19PshjkKZFKmiYa8yyp1u4zUDs
vbnjoobVooou8eoJPenp3ywkH7/jzRKv0bFpJguSPwNrmsrFbhZrECwLmhG+/CwqyRzBfmEsUSxi
tf7Wnga/5FEkNVZydCQrceF1wJGgpzzdjZ4r9u7kCrn3DThfrG1oM2wpbQAG8WGcxCi1IsEDBNdr
VeIuvK4qpTKr396MzfQ3qQMDAdc2ahtRCGBhP/S2adUNz9AblexBtrv01Pg8xfJICYHeFbyjjcSr
RatyU6VXrDpNWYpgSotTkqW6G7iEYdA5iRG4mBB3iMidGkvaB7AxnlhnpRxNWWhnt11ULdW8M+Oc
vTfJ5DaKHLCFpAgGtoE/jUOpVEb9p4QY2yzhTFyxLRUhA2t38XvPfdt6DtHRS/KFrvUgb98fYBDS
PGn2l/Nb+BOljYyQV5+N3Y/Oe6nyku0j37RRRUz3QynjFi84bUCzj+Ys40o0Yqq/HAJ4gxkMylRL
V6LBHNn5iQwHxww/IgZXM6ShtClKShLOL8RpyruEMfU5MJDRw0oq1FYEM5oU5xuMp8L0sI6EMNCX
Cg4WFsvYcTAE8HNsKgSIcNt+kpKK1xEobXxZTlbZtb1v/cMaCmzGu0pRlJzwFiqgQDiSHvr2CdGq
LN1tgcQHKlsiTrP/IzMiEo1pBxzQrTIy/mtXED9t8QaGDLZZGGDGlsSmtBewz4IMfb8KFFu6f7+P
FyEIiMzAwYGQr21KpadlbS4q37A1gAT3rF0V9OUkP0Q9tyXlxNYsyK7iBagYKVhf0jTw49UhSKU8
pqhbQvkag01DkOuhzL2mRyJXUxfZBPYPGLv1a7sgXoalPJ2uUxPSGasPuMX2SD9PSxqLLhg1f+sD
jP4J4ALJkRdp5rq7ZqhtEj3LQgScHQ+7vOZkYq22EoAM5e34fINs/dii+MNYkdywL5LVZEM9QkNV
LM162VG4dfktdvxySCkCv3Q1FnPcRxTYqrARchnUk+xSeuyOYncMuxbnWATWptWwwN2NMo8o8Jd5
e9MQglvQ/MSvy668FbYOkCQdKDP3OAQzEKR+Lfe6EevQxe3FuBPmDZfUbeKV5IoXvTwhc+ajUUuN
I4XbRoq2X37zU66mWeogf9ZTKrt6Knqhw0vuo3uiWAdTJxBAb5W6y9Ebo+J8PMwZXQ8IMydWMc20
eysRqOE+uG0qPunMtM10KgixhDOv0htrm83lnFnXtUp1Z79yi6s5EZPhG8EFNUbLrUKREzYHBZhF
+ZUDQzSBo/2lqsWerZQ+v9LY6ClR1ZHc64qnvRbctOCHe8IfAD8k3DtECIZv/6TJWSAUoLwsxb3G
haAhqtmTypZkE0HZgKzIq27+cfL+kYW1ZrBG3FXp95YX8osxz0n3YG+MZSY874abIEkd4ra1B7lK
rn7h1Q+IGPwb+xjPy77qck2tTOFCOraxQNSSpiKIQCLkj/8o136WNDiY6J3nOyWJl3D5SITFBYh5
n7dSLAqraw4NzQxPB9rpZaZ8J7T8SuDHoOM/9kG9t9EReso5xt/A893fJv/46R33RQNC01bwp2EF
4Dt0ZhqUK3LZmtzjye/o4SyU6HYqQE0YdmrfjO8NsZgTLJoSUy8hDgwldNKagDgo7q0zo5YygknJ
7C6YHtATVb6It+Wqsf+W6kHCyITvLIPHUMGQnZlWrCyjTNbzwdEkjZ3EudH0+Wz1tiPpIG6wYpMY
u0WQsg9iGsNWSbaNSrHzyhoBXjdIhEgNGDxrfnyuTv47HK99Fb01dtHB5YHOFStLu2CSQvoIlQkx
ilJSe9SM4dbgmzAWcpGmHoC+3IAZCy99JuC7dTcDxhvkfcwiyZtt3yuTjqIRDxLoKgvpyfRvihUB
YLPGu8yrfW647S26pkSTDcyrXE5zbpsoYBW88k7gTgbVDLGO6xUmmIh/dKgIHRUYSjA9ZNtXWhgF
Jy0W3z+uH98qSUcSADzLetKv/dd2N/L2BsHmxefL40YaI4IuudpJiP/smf1GF8jx7dwgAjttfC9A
sl1YqqJ2GzzivhepkQ76cGdVTYWvh0dxWbBEeb3d/PDxE18MXww2nnYGwc3ITLW2nkyjVzDUxffm
DxlVlKAWycpmSuNNAXhjipROWsIYp9/g3lV/0L0ytUAL0B40SJ3MtrqPIKZrygiE4TAqCYuVRRa6
dUQf52Fa4JxvaHcfAu/ZaJeWnWTHwJrAiG6jhuBP5j6vQx8/E/eCW+KGKNFgzZDMOod4HeuuT6mC
9JnMnSFH45bUIcrZFXcDTz0V+Rnfe4lbYERuObtDVZbVBAnsSAtiXRQZgMyuXAaE7VQ25abow++D
vv8COEoyZw+5yrTUrfALB4NMAJBjP09NZJfeadosl+kDEgUqZV4+6kpfviYAK0HBFZMqdpzjPq9r
jsiPSGWuY+4eKBtqCYiqpmMiS+lU92mrNsMFLJRgpgXn2C03zTijndaTyX7LHcdddhvQ3nkGd0gl
vyv2mat2dP9V/8mrQcw0lzS/vw73RJkAOeFJ22LcSTHffINTlB0NBvY7Cqfeve6dxBbZEdWQ6VpW
1RUziGEdhRJAg97l/t4Eb7sCznV6pIuxBTvdqn6GVLtFlaRoMXwi+qxgEc8l+U54OXickhEKlp/H
Jh5fIKNjOy6uBe53zLHIh+cRSUXlbGy2IZL1pC5I16AGywzg4eh+jzhSCf9PyRaWkytZo5cQ+NJa
KWAYQDGltspwjBpS/5hMgRlgPSBwtCpOC8QHBqDbFf22L7Z3fG3sibz1Y/TROTkL1kkXMquYyeuC
iQI7DQoMP/ex9K6yYkladvLfw+S+OjQo4w8Svp1k281vRzGWWMuY6NpXrvKhDvJGNm4CSFL17uvL
5ZHcTHmCAOJzwNVskB7GaUPmfZJX0WY3ivfzcrwv2hMWYio7KE93LBAkS/4S5Z1ixe0QBHUUJalk
diUf/vTe+gKqazeDqaYTcw54MsboSBVvd2a7oZpCXW0X1QY8bSnVhQcUkAcsuqM6Sody8BiK/wwj
ZbpKRBwFr/KmzP2fQzv1xK/T0YYt+c4EL46u4maKmP5ZWdNzRsZdsgwPtpEXYu/VLqB33bgMoQa9
mPOYdj6Vc7T9/2zuyfMXDp/8u8b2M+t8QMtYg5ipKSH+/AbbFb+RgxIj0oAAfAPNJ5fH6WHL56gJ
qYQIkDOAiARWyrl5NI3iZO4vzXQ8Eg+80klhAbSOtVj/yuWn6wr93j5rqxmE4FjjdtSuGjZpwXTA
93HqXz1EzZrNdUBvLjdJIvRNZXc78o1nK1g/nDq6OahyuOdd4kVhdvPps5yXqImpnXUY0np+/4FR
87FO6a4R7WGSGlS2QK2IEDe0sGoQ/qNOn9DrzxWnodLISUl9kNMtPrzxTosK6Mr3zdXAmt//gtlk
xjxVI9AZK2kfjxW46TowIPfKj1e/hexb/B0x33cUaG4lFoNYiNUFdTLJwkpaBK8/k2sLj8uy+zhl
iKx/V0SnZcqjjfJOgQLQaaZsXlmm6rZs1xd2ZcRKtUhdpfnNKoIw0A7NMheY+hL2eyxgn1Ipeajf
v+jx/u9d5NXkfY352zxHgjUUVv4oKbh9Qy9mXtnabG6MQi1O5Mg6WLvpuyV8GFgGBWOnuwxm+JJ7
3hdCEt/YqfMyxuvBZB8FoomAPAWI0I8rVnMrvVDVTq5R8woQlbJY0VfcjYfYLy9TQT74/Xzh+0jq
Xldmfq9PkGJy81Ctd+hQu+uQ1Xd4hY0r4+xfXDOvcGb7Ncq6AW3rbvYKPpovU1BOH1vomRh1qC9L
1xDTSs0HxvxYrywwuObHDrcc7dXybVAh9MQFz/o6gpImcguv7G3N9wT0Z9ENpC4sBvJ8/HHEKkdd
TjWKMVTC9y9XZX99zc+u92tVLnxNeTOxuC0OxVrG0tBzaQxAd5A7wOu/VbvHZW+0f1Hd/rkZa5tX
2WAbf7YU4IF+nrNg+3rBDs4WFsMBKKmpObFvDXefEUrl2ypxZC5/9S8fE6T4JtK6m8DA7c9J7xO0
enqVVbVCMyOOgYaAMJcQKbK9oXYNPOmR6JybUuQiEJA6+KLPBbO9e4lDSy/aaHJAUBYc7j4YgzfR
XZuQ1nbW95KJHP8tZWIi1SlpAtkmBDRxsgHoYrbxF9049xi64Pf0Zawde6lNhF/mPMgkn4jYGm8a
Xy9IsGDTXQGLGWVgTlwp9y5IOVnqq3P3mBAsG8mCXk1IbdbbAj+0feldD/tIr8P6esY9l0tMksjX
iqxwkrEKrjcnZh9rkYpSh5Llzmwe2PPTAzuSrNjiBNoP93yxMKEsmTOmVIYplpsx2DXmwDeVjSqh
FdhT9fuIz/j+bFoz3W/HvYfUJRnfy2pFfEMMIf886HNcxvyYFm5s6F9wvL5bxzARrsluoMdCXHjr
oo41N4J/BdVhxSRQD5epxYXrToFBJGTMLicuyKL6bnJEXNymzQYX+VcsphVc1ZJKv0NWjJ0yJizo
XLDv6FxNdL/tUMwSFjnii4PqXUJkOw68vSUxq+iKHh8zNsE19MaUU67whcevDRYNoUdlaoxOQNUC
wtPKo4ZS6uEj0rmwcZSfvG5b9wDvHRoAMZkanWMrPgXTVAJogZTuFAc5wEuy/JvuHBiaR0TT9Uuf
ZOBKCxTu/abuNDCVOs7togVOwmoTahRfTVILN4K91SbmSvOgxDxmG/U1n3Adr61+MjxiRcEGDShK
cMoSj+IDJ26jetCniB+dKT5cGp8Qz+txDFvADMqU5v7w06eimw3begkwn7duDlU+SBVXu4lBHMrO
Lx+hCcdtzNc+tSKbSiHJCBY2SMTzHP2Zdt1kCqDL02DXi7Km1Nwdx35eZiJ4uYzcMfOSniXMr6SB
svEwJ5mes8dMl3lBHHXcErCtWciDR8ifD1oyODT8hSFG9EIDMoO3unZ6vaUO4uflWog7oKQsaTcb
8fqH747BIilLMYdiVWaosSrONf96dq6Ck5VswEJeGd+gXryYfIdRIxmsO6AxwmUlLteys1svBaEl
NnkTzk7WIFIpXV30dDXlYtE1awLUK5+gnP9B4wQxF2SLeJ3MtfGmLuSJL6iJ8oxFIZ5uDI2j5ba5
kWUd3amFJfzOJPckPjpXwbxYlND4jbCgL6i9aCAPDcRtkMhxHnJdtrMkO9M36K7o8Ifm5eD53VT4
83fpgpTS3A3wFuZNsIBUgdYnX6C2DFm6zNuVeTL5G4vAVl2hnvWEBLocDczz1HwXfMlVzTORyjW/
ywJq6PDhtlGCgLxIZojj/xXOwOHt3rmAZWFJwIobuSkxGeQLGyGLhB3pvxtfgAG8rxVSFT2vUILm
v1mx/nu+I1jRR14WB/nuocyFFpA15Kl9XciFI1OkDRD5O5zNTuv9+udRNpTGWghWhODalkm/2kL6
AS4rhlKb3yuNw0iWy9xbINXfwqDwm8bdXIPRYM9sV29irUOatAPN0ThIrsFaBRyL1N2lXaJ5Uifj
Va66GrHqFTbpAG0X+jTGsUkmO62Z58JSjSIHPwchFai/Ktkxnue8IDi/HDITm6noLFwgyLXboZVK
QYEMGeq2tn4T5/niIBjxrig2VW2PfZ+Kbf8+f3rhvKmd0FQMLxR4+m3DaqKRh9u6Pp4MQAOrAjJu
nCSwsSddOX28DPvh9d2Tss8WKKf4qtJXyDXuOL4HfcaDBhrJOedkqmBem/C5eTHEXgloZgy4E8V3
mmC0/YBxga9jnudpiaH9SsHn4vkttCnCx2Tzfwxr0URglKBrkVgC3q9W46jfucnkHz6yTQG38Gpp
jad9A4kxC5ntqvii+SoGadI6zivbW//nqxobEsanWqtbV+iRZ/96JB/bmhV7KKgY/8aVg4XRatWz
Q92CocZFnCXVzA2oZtd15uNIlozXPzdFkXbmXzWmCLgVCp/7jY0wIrkCw6kviE1s4NimM3slapeg
nOFqXbwUE1b0qwLCAjS3smbjOgvigWu58+bqMO4e6DDcecDMrCE3qjLtzNCFoCA1IEPMorJ6ReL2
e0RipdTBIiME6XDgV5E7jmXWtnwp5RCPzQgVzvazdagny1Oy/QNLgp5kcBwS9IMUBRiO2diK+VAm
vpGicQ1Dqe+wcW1mg/XFGcEEYMfMU4cwa/ZBjjUigkOVQrHX5OQ3608wYFBdSsd9JK2De/ZoXAAn
4CRygxZBuBEvVuRQ0GHHoMj+yvy5XfctO+l9VIe8AWwqUKygQ3Vp+qpIEKf7bNA6cMCG+FkZHbRp
q8FPrq85ozMVDAWwN7oHzWkzKEPhtGcw8HIq4qMudc+8iG5p1bfmFo/Di3Lsow3kjp/AaNmIbBAb
a3Mm9wIC0pLwsfDBVvHhqWu82em/VHUgGbV8r4k7uvm3ADFwCl1Y+w8NLBb47uXL6mf/dBaUZGpZ
L8pgddkE+Fkm82KWYQ4HcINOHzj17RBmmsZqiS2QAbMOwh+gu9YehtRseCPWYmjMED72srPEB3Ej
q9cJ6q5Y2mKeO/kxGEXZ1nESZMKmkmpqYtQToFAKlt1uDlXyFwO7XTC84be4m/6k3SwuXCD6bbFs
Hauq1G3oE5xS8J3CDO9n4M5KOxPLYvB8eCyzig0iX7eL0ZRh7G1BNoidsnN/ep6IJp94eWldYOF2
Jtxjmw63UE+AcVSFnJeVe8/0hdYWRXICNt8LcQMgjz7Luw8TjqyP4wyzBLu1yJ98SaGeEfTVIpC8
1Sk0FJ0SkqPsuTialnVTO8/SU0Tvbl4+EG+fzrllk7FbFmmN2+R4w2XNPzgXod5BG9fvWowUPdoq
a+O990R9Ma4hOnNGsFzI1eiulbG2R2vuSwS96nSNd2O8RIJLEEEyyNhlfl2oBXZdtYSmUWPMTafi
9JNk3upn6ndBEaiErbriuo3k/sm6BfY8k3WXLFo81va04I/qJr/jgzdebKG1vtmT6BLAO55C7hyz
Dp6qdAHsgBkZFLN49Hoz3eQPv7Ys3+DXLeKONiDhTtRR2ObWGj+pmUZ+YGOiyDYXb9yTFC90hVgp
LzIJXD7FUvvAV2jczwzAY33TNVbkZGERjI2tcSDCZCHLpHL73/jEkJMj9ObwPHhATpEWqkv7FGPH
12VQlzBm2I4aCM21f7UWGKY7GSauWGwpOo6gse75f6Al0njr5wk+foJEXXhIRn7jCXxvIgGJg+an
vQWyQPvI3D5XEZrNSBfrYdt+3GrRXiVrfeDAoa65GCUZJfcrx2CAtMTVJZ78Knh8nt+2Xo3WFMax
vQ/1M1BCN5RmLeo8dW+yXwIfQwwzZgJdBiliw/Yipo2vc+/17BhDz9rCoeYdq9jLCn6VshlNT69b
xG1AItZA3MfxeXwNta6B4SpcHKr37O+LcOFDueOsKbAQJJ1Cr/eywUSrILEuqqAr061ardq2D/it
rEnKyC0ZpNJHOtpg6NTYBFaztX2cLKNOSyPPY76jcoiNQoQ0Dw0yLCBqIgKZ/yD3qrlO3LZdiICa
ps+8xX1a2HlT0BB2/B9d1F98oez+XLRu+aNjVis6/Snu2R5swqVh1EXNXTYuTjoby+AYsMBT83y8
iqvE0is36TDjs0es11kAN2BHO+5KU4WEafXNEsol2jCe6foLOvQOB/TAdxfWZ0pwTwNb9nuiQUnN
diAdQQT3DPOCOkRlEeMPeoMx0t8cx7Dqc2nNCemYYeaRbF4iWny0D9DSCQd9L1qEHIyV7vugfrMO
f9kdPFefqL8UJiVLDojq5mgXA1OLLaa4wWFq+I0i5qoCCPwdwkNVbANw4Gn9seNxZ4kYZkDO9DeB
uthZuCtdv5jD5ZYBqd00mTfo+ld0w6QQSiv+7aWUzD46XMf7V8Wjxcvftt/I3Fm7bhrbJjFxkF8j
4w9uQS5BGJTn5HOLcZ2jhD4Yxafu+ofpAD0lVu16N/teFIA1KKWpmfmGDwNlcebQpKyEhGBs5AKD
i2LmIygG+YPhQGUgir04H/riOOhGAjpEzVKa2jJG1Xy/6nJUsxaXQ/IL4Sy3mAspQh3+MFb3lvLp
pT3b3MorboZBNP4bNxqqn0874XoI1y5SINZols93guuquPvpge+o/Jpza7zgrYQfu3XEn7rfyFsm
zJZBEUOzAImJqU2BD+gFuhihAF0M5jV+lyl20fPzt0FP1uIcGoo2OrJk10kkFkr3gPeAhw6SIzfp
+DfS/LQmyMg8d+kiD7wz7n/t9m0pCAy5HNCyRnFhN2oC6WfeDP5wdPv7nSmjCR/Mj4VYSJcdWXDu
Cul27z3TBPcRudsVv495vp6mgXLAKkF4Y0YEncIj6JR0yKBhzDEHFRPkou2QfdYsopDiiIM3CB/Z
9mFf1rM7nwRMKA3777G45WfU1kLXSxjVt9GNDm0SWHWmOa4Eu9zcruGZ3hAsDur5cmDk2b6bvLoP
gHawTt+Ld+ygG2zdHHCPXaaPjOBDk5FSHLEzUtFPpDJQCTBPbLNIkJGLOr7FWHKnNB8vzhDyb7nU
RO+zKnPCNQTOdUjOfSu6YSoe8WPHwXv5Ge9jKdO44SYabPC/1nDD0ka0a4XKdsrhMfH8vVgkyQch
9f1ULee6asvy7bSlfDhSbXU1VRRwyhB6dApFqz86PBy4WBMhLP4rgRPrNNbe453PmuSo/n2nsD70
Yw0MGWJgTyE/CJD+I7cs+lnAcm5r1j0wfjXGqELfMymckRC7lpkALvl3NdRkRmO7Ch6b7H6LjqUG
vyVngB2nncy/pI4sokvlIRycHugqpGbnHVy+pUWMf27SclX551hae2lZCW84diDWBOPT66rwkexp
dZFliNX79pJ+7VqjdNZFe+1JbCEdV2HJYlBlde2V9a9oV47VyFQVAKr2mFdyMMtWcXrxeV81DfF5
Qo3+QkD5ayQX95pHlHSYZfeqbG6n6+8F4sEP/XFM2o2EzE0kpaJXLeIVAgQ/NzH5xUJ/yOkTTVx8
jY9BtFD8ITeHDExQWjIP5eaMr4z4J5G7axJb0gt/KUFHsoQabNWMuC6SjImLRdmlPPsroRWqb17o
wOfT4cc1LB5iF488vByV2iQkKKZwYevgBNy91+VoKswbx6erGKKQC2jKIwSXY4Y7s+nvP07x52ho
aDDcOs27Z0alEBAlUevCZ5JTYGs5Pw2Chd6RUmV4HkCRhamDK/qkAHehB7b7kgO9gx6cQENhPxY3
z9N1X0TyVIdQaWZOWVXO7vRFaTLClp3HIwZCR8OOUEjkzzEuypcF7l6zMarK/MsP+GOECffwIq6o
2pZdqNdioX4BIyA5wBBLPM6oz0KaweS8CRUKpOqjIViHSuc/Txdio11pitnTgQQ1ohqULrWUebiL
69rXg3uL9jgw3lCxmorgcQwO+srUEkPE9WBbEYqnzEoOB0CudhOrVeZjDsPNjlxlHcwtTr7XoZlX
I6JX/OkPjguNvL3iRmGgoW/ceedvc07tgqn1BybeRsMRW0k/ZP+YeN5Zc3qM2NI3/BPL8Y4xifpg
jPUEt4kJ9ugcOEMYlt82wuHk2s9af/+JqMEoChtW7qUYyURUH9t0BRMTZC6g2nGECJaWVHJ2rYDY
mwok1QEpWo8TY/ru6gjw6JTEv0KQfMzfL6qcCM8RtLsCGBcFaFx+IqdvJgYGDljc6vCatEue0zuA
5kiHCHHka8mZZtjHv7sAYM72e2IXvQOmz4zuSe0R4wrWfZgq4aqDiokWcgyV0MxgXjPBeusddzVt
elBlPPbbJSMFAmvWEWZ89VDldXnLtGz3dw4GzzXaLZRPlUYXFrpUteMxZd85731EzdNNpohs1Rpk
F2ANqzeoD3t07WEzUqljmv/9GFplpRTAVIe+GZCGTwN30kxW/0iLfYVNRNtryvHUWud/SdTKeb6l
eb9CnW9L+k7b2c3plMEJNhe6ZIbob2zPIw1cKvoEZUtSjvBdnZvPLsHq47/FeyKWHRePbLB10IM3
cJliYVFkmaI2icByYMyqYfDryqRwmg2fyeSnEUqTs7i9iUvcOUtgZ8nOF+kwI6tYNuHvEnwXYAwD
3ApiFnvSIrXrk+9zvNbLSA+KSdnKUTFzisd86BGcZj95+vdLh+kndqJjA0DBMj5cJUVBBWy4uNDn
7s9BbsP+GYJuiAnsEqdZ3UEinpSAboTCM3KlCFtx6GL7kZgOhB1QIVm4+nIq2r9ndVoNjPkKAmB0
zTTXa5B6x9ad7PF288aM/5sAYhKvV7aOfRQ/yeNN697cdVXHXIYuJ/0YFZ+onVPRthf03nDnaH0j
hAYDrAHBj3wntk5qYkfcvWXtHRc9A3yzqGtr6TRBkVP9wsNuTbba4GEldPvuqh8ZiEuVrBLdEASY
U1sxseCGydcZqzyj3SRC41OMY/Ki8+SlK+Jk1BADalYQcg6eFjzDnZzMcEnsLmS95f/y2vQjxVTB
2JN4I2Tz2bI3dSgFV2hnF2ygu9AlWYomdDagdhZZvTJonTHVK8y+iX2X5ZK+ysDhcTo9KuC6lzhT
wJEoWn8zwMpYpJPtRqG7MbTnBf5kw9xKJXzmwkg3q2ittojAZVs+FAj4V5kqjoKSnGtnorynfCKU
U+O0H3GQpKev1bbpfQnBpOUC6JSwmL7VWkg80RChbCvnUlObtMai9yZ90POMWXEQPlEsS/Ei+Fyz
QQgiLzrBmIh9z4OlTeHkjZ6rM1TIYswmBTYOoZ80IBtlzz7sF/RSN8d3B6XNwMpn3JrnfZXiJbRp
GD8/5Dkcq/+gsealYDR/wTy4kwV+qhdSYKAhYL92ZJPhYf1MmriRSLS3+PzeXQMGROOxuJ/4VnbP
p1FZ4hl8DvaS3hkifD78Bz/0Zup2isv0KUjgJWzI0r53g8DuYk4RRHlHnYu1qtYJkiW8ZTpkw+Af
nAgN/hS7lVG4mLlOnqVg6jSnd/51rbk6VpGBFcLtoaAax7+P++isUrp6vWPvPkC6kxUOw7E3X9P3
68+96KPnWpJV38JW7AnB9zoaDQn/GC11kqc3KFdAmkk56zhdey1zhNfXYGKlZscr/293NxH+rRRz
34SgQRexULcM/QETmgM5NaxDMs6LB0DuioJnWu+ooGO8+UfpsGrIbhrXPzOPWnloWpYHt60YmdKy
I5eWzBLei2+rGKmNMIKzRsfEUo9PkdStlqyNa8UiDFqfGY2HS1msfTCZksiT21vOPFqQOt3hZkCM
pFUy5fbU6NxI3TgAXzGq/Ja3+6tS1e1gvwpGDXebBA6dUYkK9yu2YHcXh011GEVcPBtdZNtre/TZ
GbPITqz00pupEyilz9caUu4WczEw2z3NiYD1uzwXnLK4fVwHsGXDaSyOzGZ1WivMcbOFpcqsybB2
t7Ri8Oo2FYrxysOtDcL0hlKl9zJKtZEtba+WYyf4ffYk/8G3T+ihy60PizWWwTZJQAjkY5hQ8Ptd
ZnnnPBXVIW+Ip8YhVWCKlgskPDIHzhv4inLdaI3tFV3rf8oxpVFyQlyqVMbntJlJcvAFgucEefug
IePnxuD0icKaoqSvHZCCgjJ6Z0Nb4WG3IClb23b41ZK2eH5gkcjGl9ygWJRuuXksD2c7ONNI3u2e
mRPNo4DoR47w/+DHjqAgCuEUsrFRCsUkTKV+/1kx6T9PDFVlRaJ0J+cPN1KQ4R4PUyE2q72ln9S1
n0D/AWNbBEet4lrwBU6KkeiAHAnJpfcLLbI2thcireYZmNmkrsVKp4EfCYW0OgD0agr4G4WwkhL5
zjfQnVLAJqi2JElK/7ocjammVKxzFSXzYguOaAMHhYAqt81ghdHUbKd+ajfdkrv99o0Ku+dbHCMp
/bUagSLHQ0m9nINXrio+r6HmcqRo/JNUqiBrwNQcBdi4W+PBoSt9f3TyUbcUZiNUWWbFIU4phXag
zZJSku761p5CoSlnThA9MCPOSXpLGIm1Jl7qczPwTQ1dUEnGweHLbEGI6wJYQezBj4Wa6+sBKEjT
yizzgRt+l3CRTjFscqZTxsgvJr1oUOstKfGBIqpBD4ic8qG44Dhs9Y8KK2+dBsksmDX/Gvd32CDP
7YHQW2t2c86FhNU+zD99oQo71oRQb01N4AKFLcpHKZhNGjU17zE0/LNGj6NtxafpPRIYJ7OKLc03
lzSXMTtoAxMLCabiK4XfD5Ee1ATdw631eRj94smzJvWFg/D8NBDNvOiS3CuC4gzbAvlV+muoxrqG
R3RmnzyHey32EEwUUgFZM7o9sChhySeRw9U7cLIUJs1thiilRaNVhQs+36AhyB8YTW035JKiJc03
MfN3r/fy4Xnn2K8YSleRdCDojuV3myE5cLXs6VfTuPe4YEK9gqsL17hARzDXCed8yz0M99HJ24lb
LXflyIxCNSwHS3sJ5TXsc1a41OfbMy6jjRkJkkn3xi7QVhLIIMYjhuo5n7tkQ4tA9xHkpvlGm4pS
Nabqre+KWplNlxBqU+KX9QI8nqIPuzqsS8HtxnzAG2yMK5Q2ni4uarsHA4J+/QmQ4x8to5eTKwer
2T3DagSWyVpgzfdDoxehEZdIYkDtXpA/WuGFBwVtK83Q2SLE65ZVwRG7D7skSLXugfLFtkzPf5u+
XrWQtHLvU/79WoYzBN1liEAIolP2Hl1+dfUcvSTsgXdcw1djP+qwaC8TbCdPFZo7JzPRKCH2kpXD
uR0ZubgJbXwi9h0zDYrGui3Q4uodTxS446NbMwC8dRfUy3QJaVU5diNKSKTc+GQ6s0Nl4AKWM6bL
hUKNBi09MXxMBFTg3Mj/hus0/NuZ04Oitds7QnhuC0OXqXDiQX8dhlAbHp4PwpfavnQWWj/TQbc7
P3G3alK780fIYVqvU7b+bNtRaOp2aS/ZexjwD+9WZG3CfPUqb+/5hOIkSvEVN60ZocXeBYp7qzZ5
5UYLefIVaUD/DCXB13PRI4LWt1eINjDUXhcU9wvnl8XJbTrUw8OW/8NjmuPgy54V3EUEiICFDMVk
J9M+Hls+VF2vQ8z+JS9YezxRDR8qRgu3z24bMEhCiujGLweIZkYrpW+KO7Ot62mT58hV3hB5mJYY
QVoXFcakKN+n0kRAu2on2xXvEtYsHWDBRETW5YPnzaqSb3kESdwbxT3+AtwejkpV+Pc+7CgIFURI
iOefJYpQ2jdjeiNqBQMN0Wko0pqHu/mqVGSw3IHe2zi9SrKzxwZOKAzynTYL1J7yx6/f1BC338xD
sWiSqyd5lTdzJxv0vpECc9CpormzPZzw9KdWxKXYgBxxb/5O3HPQFHQQtlJBhITUgQGycm00iwvw
Ej+aaDhPfrDnr0YDL6nlLYEz9qH3+HERDueE/xK5akjveLZ2LsP0xWEt+wjZcdbZUCBAiWrGOBoY
rXOLVL9mCpogR72zQa8i9VhzpUi0sfl5GqwDFj2zL6g10/KOjO4WqNo5NeOCvwe3Bhv69q6TcMJe
qTuI1yIkUI8ieG0bVc8AkwJokVahqNZEFL4+3gh4rqaKwMyIlcLh/5jHzXK+tiZHsORbtG2B5nNP
I53VOiKR0Psk/6Z6hBGBR8RjKeLfzK4UeUNedZiOW5LjQiFTopP0+7WsECsrP+1JyveTA8jQQ2QZ
LrxbsTmbF2zZ1P/hl7by/3+w4LSFLtAEoFDOeZhbHgwdGgg/5jVzTZpRSjeKx52IQXlObi6pmiiS
3631mmYIu4J/whQ66Nr9ZoC/oQEEjpwu3cxgHLlPigCRmE8o4sztgprrPoOEr1lf4ORoQmatnaKG
ZOS+YSNGWhGvle7zPW68+ox7AmYARM//vXJKMgUN+6Si0/uYOzCb6foZOesxOPxRNM8kI4yngtZK
EZUuNn1Rci8fNe1aF/JgzlVIj5F+42wLGRCAyyCGNbY7qk7T4AntS/3+/chKcWA7SDwz1FOxI+Jn
I41DY2VFyQsmVuAf4wwnupnH5TCaaEBe8TDGU308BBrACT2CiD0Ex4MdyhnGuxE7Q55nhMDhKK+j
o/fDnVRzJS76GySM9RcwZi6yV7Hs4EgpgoA3SpWZDYOvMmRePi59RZWe5c6NAHV+tW8FEv0sxQax
i87x+JJo3zdw3tIoBv9bXFCny4LH5AhtXTiDQnfsVtSuTxe4erOY53cDOMB0zabHWe2KVnAQNrpV
xMbBqmaOiPBtGi5BLyQ2+/7jROwS5eHo0ARuVUXZd5QfRLJH4udafiPxlGswXx7rBLc2rNwvD2eH
byGRqYGgS+w7gVLRnzM/X6VzdCHJhGWsY72Gzv5kiODaPXdClSIiN4DrZPh1xE3EmWQS/6S4d6z6
TT+SWH+dnCk+L/RyBC8gg0cvCtajlei3WNVZsX09Vw6fCK898S7gMs24PPwg6fi16kzxzhqusM81
2hLTjhxMCeP2SnjeCQaC2g37Qw6RpU9oSG9hrNyZVGmXzh4+FruM6GOLo+//rN7jmHSq0S/Ad0xG
8PeHTZgQHBNdyoaEkH7oe3QC8v6nXjZKpKSQLAlDORigZ553vM1NcGuIQSYKugqx8iyDkQQ4tL8g
AzvuJWWUB7wCFsZYn3EuUC08cg4leVpx5WBkq2nKmcZNqpx+6xYT3AZbSPn4Xyg5WcmsqNR9GYS7
J/nkt5EXKxetmk5n82CveGBEo2Z+vhUDF3v9BHBxyUpM3K5ZO3CRNxcnce/T1WftE5jnqpWmdHjg
Y2goyVj5Eb624ouKYCxQHZ8eSX81fkFj1ireFnKzqirMRrTArT2c9mmAm4ExjsFXMuk1+6mwH6yi
XEv52mTSCLcWnSmwSXNPJSbLj0BwEDzpYHZ0ksTCXepEJwOkNoDxkGRCWzE6ZeZd45jSDxDzEMNt
U8nxmtbBBx3E8WdsGMtm/yMgL3k24jn74XDNFl8Bs5HfcgODW5TuG1O8abF56+oukdU3P9oCRB34
6Y8616DoXiGC5hyvkQupQeZadVyQeNWY9EyIcpQFV7lxTzaw7g2qAz4blyk5vZ4iXMJXiXoDU7oe
Nz3+hRM0FW0I5UMr60vAu0ege8o01cBQ/TohGhD4s5GMtfx0yGECRfbjPsnSUtqOFGb1jlIIonFz
/TiMsXHDqfmptQmR825rK9GmmhXo9iPiBbii5QFrybVkiDGNVXo2i+e6ACIoVU5KWVrGyJ7SwgBL
8Y2jt6WSVJ+IVaoX49vvg284DrgdDPDbwRkZp0pa61duFrgT/bbLAh6oHA4esPLnmw/uWFwu9gDm
dXn5L031zIIoWh78ds4Yt/dm8l5CKqONwUA1X/3JEu0MeI/y7RR4SP7Bxxty/BPYXcwG5fHolVws
CA/6FBDRa/ipV0NLTY4Njxmm7UX53csB74v2RzOc8+vgIoJYlqATGRiau9QeRXODOa8zo5RHTafD
QdfZoiwx6/kgQGEi1Xnvg75SoJYLllMtLt3+Ns3ZA+m8J9BKgkCeyZwgP31y7RQ4Pc4hakdLrLqf
J02D4IOaAmXk5SXjiGz6LaNJsraU5UysXxn8BgX1DE8k/vRCOQoY2aQaBcz8GxXT+hl9ur0JHAmA
MREVktiUsA3ntC0WHiMQw7vMsMPEvIDUhtROQpvQZDyzFqCiS1AhDlHd0mkRf2HjGmPTlYJPB34W
KHVaiL/VQx6M8UIBed1uj2K4DrfguAzAL7cwyD47Wq132WjHzt6vfoaGQwxBoGA1PPbL/m/8P6mo
RzR8xhIrRYwC3MvaXZZ3qHdk+T9vJXRC3fXUunB4zzkQ6xEnBs01ogf/Mo/pH+PtZhuNlmwsEUX6
4LTzjiZ6s5opRpIrQQp88vQYVJuGOBvWKDg/+7PwUwEom8dZKGBseifIZ2sWsSZT0zBiJbJX2PUD
NuOVR8OErpjH61YlS68Al3Gnr0XpWZITlJzv1iz0BOBValA6a/bWFKQAtXyqpTEEPu6LeguvaCkV
H1H/LbNPg4VyPljzyAKQZlf+Tfn5DxuQJpQzYlg7MQxcaxagntXMTeoQ4026vqLCBTk3E+Bv8IjF
STfpOLyI+u2Gl5/fll61rObGbgeny9OkBtDiCW7WdWOq/AM/6Es5qMHWmkZ6L7vVllnoorAHGf2j
5QypszhjSvgzlclM66t0Bs1ZK2UIWsqOGDpYbW9vTT05gcGayl7pCmJiOKDjHa9iOkOE0YsNyU8u
aIqNiLd3MTi8xlzFk8ho2IF4ke3CrYsSqVI+F0/9a4Tjwv+MfwzD5yEQPbQZyYP7e7ZDA3fiyhjE
Eg8OAJn13oB7V6ODwL1v00eiRtM07tKfifAgHvpNFlgbaUoaMJFFloIVy8zQh0sRpnUwto8MV+Pd
k7kRXTNmYV2DS3b7ti456zyoQGjyF4GvA3bBH0zBFUlVNet8M4AhKIfnyh/G86sOOZ+2gmEJSm6m
aH8s+8wDtNWiRqaZlVW1Sf6la/6rGO6OV8ZLiSOd2U72W1BDUwSeL9MnDhUzlNKObORriUvgbuyI
iWPtKgnEmT6mBi5sIsK3aXOcw88VFLBxpoLFHicPYg649FmXMqM2SbBvNHPI/8AtFXozmlhi34Ua
GgsshU6tTzNjrqhEFDQ+tOtDYyLAYOiA/n2+IxvfC6wkaDjbwmT8hBrHLLQRBrFRlLXk3Bovnz9K
l8Hkcknh2n7TdoXBWPKhjlh02CDAWLc5mXdhYMVxCwVEp21eHZ2M0mSRvMUZ7F6lgruZ11IA7jyF
10rX91Wmvu/j8fwlOXjKMl2tDFoVPPFfUHubkvid51TBme1vRVC/yE4EDoSMU2rZhFRvfXYdUVIJ
K8XAdGhinDpgPRCa6Tap1BjuGKMeD/jVjdSREkiZHkSSCJnHdZIqQqF/ly949DcM9QsgtBnM+NoJ
45+JHC9V/270mfrb8s2VSAcnjCNc+6wVei4Lh87DUr/Sj6mrCYn/jTe52vS6pX1GaqkWdk/Ygy/i
XPlY76RPmFSc61GjW54L9M2GwS1OhnBRYy504l1yRXHlJujecdCGy32sFWZ2f2aUgmI5E92nUu0y
Sn1RiuyoMyKxR82+1jbFfVV5+uWpN0h5ne5kHmGT4mjQkOJ19oMiLTfaW2YcY9gYlGQB/JSbmKFG
E2MD6k4ksvN55dNClHPoCxDzv1Lags6QGdoOG1F06FgDp7yxy+lgbqnqRR/hPtI25+PuZkvz3hkN
GVoHNV0RTQQP8HMreP5eTHc4oA9sPgNdoZLlOx8v2jkoFCZdH1cjPqCkacAU8eCxqJ4tduoW8EFS
gaXLOBoLfrhU/adm3CHQDpkXDDrUpW53OmtIW99ldN4H6ZSzKyxzDYlnX9edikeg3u7Gw50/zHA0
sOs6L7kEk14KRuKF50HtyzTESpTBvPykdEsy/ndKyzxxTBbiUTphz88JUQeo/k/1FZAMCxjmm1k0
qyrMHUVqPFBmIL6phqApMH7TEChHcicOXxS7JmI6PUXJeoxtVH4l3qcl7FyNjy9mYbXM37RmsKL4
APZf+8wVowj/fJZSx3qJEh2FjkYDcU8+e8uOD6UKCXzPOthNEkQZnzZakL81/G1O765Sn9U/JjyQ
l7H100YiACGudFecTSLjIRlJTsKqZTCD+WeBTndtC6F6YhDU68XyjV7XInGoizyoOgRegDl9qTGP
+RaJfN7Qc7zSzNlObpWaYkypefbShWvSs+23+toeijL+zOKttXlZiUgWdvQur/91ffzXaI4+F9Ct
ONSyiAdZTjrF0H59/MOhQNY7k+XX97hWWQisPf2NOs13YrETS2OHM6lp+Ia0hS0yb02fbWeFbCqr
wBoGkjbBM5egkVjWGFryVlEXy5PNaiVLynQLMMkKfaAck3v/6T6OR9bwIagY17m2/9+WbBZ6uxH0
CJVE8/Vmthw9tjzfYLFSHQSRqL29vJvhF/Eo4zmP+uYvNLSVKqb5Jo/3xmPlbqvZ1szfU4VRiyTH
D9IFKfZEhsgzgzT0tq7J/VLtHDQO23hWwJiB42dz3QSZJdOEaq1TtTtBBXPvai5FUaX3SoGfjiWr
Ydw3QJmQMqSXeSrVKl5E0Qse4AUS1miX3zRyO4JMSZscUffgCpvBk2QG0MkTHfwZxiU677TH2Tlq
BwCnx6OmPQ9E28+AeZ30rdeFVKpJsLpnxJw0uuEshv8i2tr9q5GmIQs0GLs5VOyqcIZVkrVIrgXu
0mOQ2UFKNdIyfrU3oLIDskhwqwjGOuhUypLYo3bPCwwJft9SabPC+1tXT8eE2aoxVxnqoyC7ON3L
YnyeIWiI7bOASnc49lYPB+/15b9fkHeSr9OBi0DvUw9YNKXXhSNb+WwXzYlrFUQdpgAQiOT96Xrz
E0S1B193q5RTW9mT4uIQy3oHmPc7aZN+CQDYEEXU0FjCa0j+yWb8KTNVT7Tv8/sQsSZK92x2RQJY
26xh7BMjP32wncaYNcjrg2NJ1FHgOzTuc9+7+F/4BXBjNkljIykKwHKQYxtCAluv9fnxbGwzRzFC
wmxJPePYo44noBMInZ3CQgSiEzLBEkuRZayWokD39CwyAC8zr3g0GCkFENwVt8NEpGYQRIdm/JSZ
IC/IOjwO3nf1e8gKTQJnTprYgvn/T7tUKTKX/7++Lmk/MwAYBGvBQldi4t6aOhaRqZfqH6H8d/A8
k+vUF49kkhdODR1QAZrfcZsApDV3AtOnKuPgWr2e2mwtDBBtHGgKbZcRQYn9cVweK0Cerm0R1IuW
3eJw1aJyBPINi2Bf4i0G8/2azLVMX9m32rgSvlOB78Hrr2BHIFiKhtedFHhfWfPfNBSRd4bTshLg
QLDrRFrMpRjk4DOr/9jI0hzdGL3sxp109KvMQMcUhu8tvL+CfD54VlaZIfi6HrKVwiWZwsYkKDiD
ZRt3loPjPWK4nr8AxS/s5/eyKgAFDA5PFYJoyVIYJTKbF7nDhg7LqU+P4Ja/kI0ljVNatImlRyLW
/LP2LQgIrU458JQ+f71tKLghnV0Ws0aFtWrW/NcrzX5V7AcCktPSfpQx2M0ZU30thZn+3WnQjOUb
MCXNMvR4HWhvBnQMWPehArUd2ufqlWXaXvMJCHkqwVwjyqOlJwqDjiWwVZtUCdQGse0awGpNc1Bo
exK7LyXDZLE5PlTmgfILaPYw514rzCReD7ZwCB1UfclEytCbhQti+So9UsrD0O9UIPzRUl89kHR9
1RDo+tVolxhylMMFSTX+1XDJP5Ekoo6Yt331S8eCwzfiiePkgEAnTZOy97f6O3Bztzr2m2Fw0U3N
/84e5y7iRYyXF8kd3szb53mjrgQyQdWLvrIprknWyJ6P8cP+bu5LWGe+Pya2fzgguEO7Qy1A8NrY
BNku0mAgAA0bhqqbjmj8vgSwXXH/HH12VQ+h5mAlT6ES5niuMtS1/Kzue0ZP3W1/YtRUm8jJrSPq
t5dw5C1MBCHfENw2/Xb5ZYCLHRF6jrt1zWDrz5EfGFP5tlyztGxyBXjUnidPnlNRCqDGMCqcAlK/
V5wh1ANTKCroNiTDr18EqaCyUAouIYMQn+l601zHqw19/kaG0N0Lomdvdf7NJxSakU0rBAiTzmp4
7hgtRpeaWwysf2K+7GRBMhjJQyelGMr9U13AjljZISQI8tpTLTPjuv5eATDgBfZS17oCcog8Wb1v
Bw2yXFv2EmDWxuZ19YCTMHRX7Ejb+h5XfCicqc96boiP8Cr6Cl5e8ybDbs5v6GwgkMISQag3tLCY
xpIWIvo92DeN6RKjHMbHXzvnYB7UnSzzqQewjVa4cmTsQA4cyD964ic/Jq1/eUQWWGy73rcMFz6f
rzC8mP+A1+PHOkD3QmUimRtN3Tcd8LJBnIwBCCU+AJo6eQ0olEkpVUUHNAn4GRcBTvfQxHl0foZg
+doIFUtfbVYmjndNcgwnaFjkwkw+T1JLLCD4bCuu+L2zBI8sl7nDbhKHDIskgBUbOQoGy4bRY9zV
3drt/40NFLqbTjEhOvfkO7KxV9FtloYP3IKi/ESfTHCkbqp5Br18tH9xFgS11FjaFmrqBgh70fG/
Vt8oAnCBQujbKtJaGr2uBrWqBTPbkBjkNwqr8ILgqwTNT41du1//ycaKmmUx5PcSPA+93SlNE5Ob
tNB0qFQaQMud3NtTtuuJjDz4Av9/hLtxhBLwuLdc1wSY6QrMFJdC7PNuSSmiLp0pBPzR2Z5C1iaR
5WqWEaOc30NAGXY6n4u+26KAftMmA6MKahfQTvrMnveIIuIjJLrlteWOUpnjRGiV+7CPs3cqtEfy
NbE0S0zMW37ezR2kmk+qiKV5Z23o7k77W80k/nPKpMOOnKnyXhha5Ab4+pT7Di9SnDYNNrzK4pwy
vvEyfUiWta3EpCMiWOL+0d143RZEiQ+qcq92sC53FaeJCA3ny+beeF/19Cr0oz82KJQmv0o6qHsR
NsGYtzWnc9cjQ7sNm8D5f1oIQHRAjtEkKvKmSljpM4CLHA3Q9+008y9OBSRBQLnI+lQIIMnaWra1
XEYY/XPTMHSwAPl89yYb9PR5U4mSdRyDaW0JrWVnwMxzi84ucBA4kgf8eIcyAAPFVCRQOEiowFlj
9p4oPUCFK/Chnzin5LJXILmicEehHw0TGltSB1sZNKw2wImmt6HknrI9oyS05y6K72MNdLpGuFiH
rE9poHic0gtsCfnahHKBvHdu9ka/oG8ARhwlnB532MqYps9Ni7dGfhRpVxC6wmf39Lhmq6eKgbK+
GbnvArkCXwYgQuRFB8ww3S1VRjZhDwn28gcne7gWNMxkntO7X5gK9Vi9/oOr13erL0nnkG+ihHpG
FurByXEA7WXjlDLBnfbbVZ95ikCe5kjAN4Ps9OVT+XNkZwXgZ3mHVj/PSlan+/YDU0N5S2Q6pAJp
6Pi+WgI/HxDMnqFejVpO8bgfcSOnUecm86/HEyJVytof3W9aJUtMldznLKZETmSMuxgz6IECXNpb
I0z8K2O4Bv302vXBpV6LfpEwWITCuw93gU1+NRjtJDddRGS2vybAYbxpf2hZb5tnBfesPBrvug0d
jd2SyjLT8admZ/G8hNQbrJsiwarF5kEyaWAjBSezoPrwykmHslNkq+HRkz42F1/+bPflS8qpaZ6/
BZmJmpPPtJub3vvmVAE+RSg3ZSY+lr6+WsFtArAmYmCaIQ+vTr9GrpX5aJWL31kyZErl7vYLFs26
oQizc58GeDMp3bfWw3Qd2TyjMHB4x1e3xxToet8+SvR8g3ZUFcAul6FYzdAGjupFeIBq3D3HAXsi
BKWCSZZ8Kv1xtUUn12UN081xraEHLh+y5VbSQ+vnOeBqoo99z/BaqUnKppXauzisgftKbvhehDKS
GNy09ws+hrp1SmLTUPKJdnqLKA7xA8cU9ElJGCpuwbjnQto0MYAwXxGEVtilUTbMoPo0CObnwSCT
hvlM2HbQ9JAhoFjUhUaF3Atd+3uhDIpXQLJ1DmIjKEN/P49V30E87ggARlLRI5ZRDuT+EvO/kzWk
OvRvVHx5RST1Gi6bQJAK9it49plE3QVDvBuRkSVyEZ7wF7G34djAEUA20sE8/Lnmn3xJZskAos5e
wvQUc2KKINIch1KwtJjcdV7tCn00ku42Ee1knpO9yStYbPbHSftBxX2fq7o/IBfgK/gXVuDRS+Jz
bYR68pToE75CxhHRUigA4+9thRhkZIVx0mN0hGNjkzNpam2jLy4vGkX2g178ftIrNNjPvGuGP3b0
CYVjaQfqi3y/LOeaQztrLHnB6Hq6/zm1Wf6jwng/7VAQ9P/zOySEG5oNP7xx+EUa2LIKU6EtLIV9
ujnkEoeLxZHa3AsKe3UxoZK4ymthlxXzPGjx6WaINGcxNG8rugUpzVdMSzuIKl7GzYjRjjMlD/F/
6rM9ZkkdSgZRwCi9N8UuB3yeelLxtusOcTn58FpkTDM0uqeBptiWRrHzF1rpB4n8jNPhcmp/eqVk
4wLfyfv13oXjGvWExYm3Mw2addwLT0lpd/C3Hvy9LDD/oLEP15GBGdGHRv1dcrSllUVfW/PNGiSi
Za4O30thCa7/JFeCH87wFnkC8Ji3Njr3BZtqn3s7K68k+FTiO8cXz5qwFbVdLEQinIb34YlugJ/p
krBGIpBRPWKBCF67uTXqOmveflPmCqMzjpVPh4tmSiEVkhXb0ez/i1P+bYg5I+gk6o744v7ellzE
6cEeCSHujINy9MXO9pDLZuuUSudEBDOtP5ImobzbD+a6VS3Ga91yToikhHPMw2pirWBtydMviPsS
VBmZAqubCUjiI3fTiZO9KH4VcC5yeCRZLiYp/Agzm0TQ0Ko53VAFkUxbnVYokwarN97e8keXd6B+
xhYEy/fqDkHn7QnIeBQeeBS8NRTayOSvbA84TD+rGs8LazT64BcTeMbL+C64NAlye3b0FE71VvFq
ONfC/BQNoHa25mFGOkXNTzA5KGlgf2iCNQgpeAcn0/sQslS5PyIyUuieb9ADmk2yPdR6S3NpLeYv
PQ724KsNn1gzKyVlOkBc7t+EJa++8ZK+BbOsjUaIAHOU642HDwuuNejhCl99NsCO/oxqxv36ewAh
YbRaETzZ47c4O67J16dX01rre38RZbS6SA+TBO9t4KDU9FFh5ZzpE6w/4GSl5Kl8EwK35EXVmKoJ
QUaHh2RXetg5XdYkZ6WGjCJUxCGStIhCjICo51OaZI0usVDS8bFcn8Pwz/uXb49QAXeXpk16k0la
3f8eE2luY7n3DpU7pJZEnBUboF54deGrYBA2bck826syKolNZQ8aN+4VQXMjoH9AtVJ3kiquw5MJ
dYyQW5VvH8IXGC1HNiFZH9qdGrfREoLzGpjIKp4iJuCL+dlM8JgRayMyrvs6lzY/+QsjmoJm+vF+
5rI23FX7ZMdFmCaeKyClvtF4+7X+GO96NTD/kAVIPoL0dBTkl/2VeiUI1ogFTZxVU0kmuTB+bsr1
TzjvkcrG+p1QwiKwiotdMAXarJTUlKg1tSYF1YPkNoVtS6EQbybe5DyJJzI58Uht0f+Nv9KqY7YV
8mrV6vkHFE+7PS5UsKN3k/Feju7vniRO05aoJ9JwBZHwCiTmAAqy3BFuj9LpMUgB9b786YB76Ady
Egs1Mw6BbPiWdrDrtLHANC5DJp1dPlUS0TYaUS4PT3s/T2JeZktjAV7CUtLqWdbMqihnSkUbmC8K
yKuzIkoLXL6BzGL56J0w6oY3ixzcxmCkLTPYiWHxI8JF6/vzUYhv2VKfo9HxkOkukNmE3DZy5y12
0YATcZmPcPD6MRV2VbKpIdJjcFJLzEz1iR22kqEFABWCWTAqcw8wvr+GMDEgtbR5D+1rmhRVGJol
nXlDJ/V242Ce+INARdlhG17wd1gH3RtKnsD3ho3RgQiXO7h/jipkjPf/15XV5S3QTTxk5SI59CS9
wEpj3+OgPHJbTtrAhm/ltTTjKLYqJNHobMfaRjXjQHYt0Zw2CdWpzF8AxxMf/G9qnkr6o9hfTXAx
UD1ruYrnBUsfw8OyEEe/b588v49obR5SkyTtKpFzC22e02by2knAvRuEazEt5jrsNB9bcmYK9erH
8gD2LbkSbS+It1ii662oUdANNJ1Pzhp3k4o2jBOCtNceGcMCIV6z/dfQJr6ZprKlqPxoCGiEjH5n
8M7pnIIeO0/KLChNSiUSaqDuenMDZZdC70a/3MS+UJ0zpPLjLNEqZ5Pz4lfqwi9JOkAV1cUbtn68
ra6Hp4WZW1x3lOZhwPr8DtY7mk++2Vk2Oks9Kfkn/agfyTqO6dQK76rEDMxrltwxk8eRbqDT5hne
32g5fqcXY9Ue+EKUTDSlvoUTrJt5l4aHe8Bv2QHqJ7XcjzGCtJ4MFNw+PltSsb14uVS78ysF68hp
Kh66JOfPWFHjnWZlAa6w1yNZophYHkXzZzr3eT/IGvYm20dzwY8fyqSONprUyfAnS4MWHLa/L9gm
xeN9+cWxbwkGsyGp8sHh+gqxYbX2Y+y6dKKgSJz+7JCbznsZDkyIgkB4YMvjuChOP0EEo4nuNcB0
KvnwouY2HIe2T4A8KBYqOgFTULSsVFsWQt2AFex8dSNocUGIO1PYrS2ZyY5dmNhg72nr+kNWJ/3g
dASgmn99uUDmR5kgAIUcjkOMZVZr1pUJpMDUyrO66d7/NppNxEjsMyGVEvcrTIJeaPSvFj/L/w7c
uYJH0zvjFJoEJDQyPElgbnPPp3atHCGuqEhmV6CdOKOfjA+zHFvu9PxBC5ZpoS1dyxd0BUr5chWU
av5imdk0cQT4Yi3OaVb6ttP6J6uwtJf6n/cIO8dJexF5W6cx/9Q5sKMc4WW5owuOJG5TaV2zU3Pb
x0046IR2rFTorpJ5H6DWhB92v9ZAzsRe8n4kmJF1Zte/pHrZcM82MlGHS02w4ErYd9org2Wq8QlM
6cByxaj/KKq9yMBFVDsKNoL9GYcpSCnUvsJ+mqmQcxPC5cTVTrKAGIwQtj5WEPWwFnT7DSyNzkIU
HYZgWWc/8OAYzjXtkKB8M3QUhZN9H3G6DIf/jEUEcCBL2bgiWDJKvVNsVeHgbQI0fBMlpRkWjgcb
UEzxP5Vf4QRN43zlYrdlkM7hLGjC0IW+3PaEMt9Oo8DI+F7ZYB2n5/i43AuL+3Aksi5o4f00pRc8
jULmjqWS4hXAcvcj9UZv4ozFvwYqWFpUmx+cu0jP5Ql9I0d6rA3wrfffl2yq3qMP1KIc/Mmwoxki
TyaAaFuellAzd0675jk/+J3xE8oXbUqtpXN2fqpGVRNCbY/cGkqc85dV8gkKiLIpEw0NxiMUw1ZB
RL8OPuKy+SRjVxRs/tRKkhRD7cYKDBSOLKrN1GI0HooHwwLcsNC21uJnFP9we7Xd4LC3jyViPTSX
UPOVH3m8FbAySKM00boAdBkUigJPOT8b9R0pcqjjkT7S2v3/A+AikMzDSboRdNFEKnNX6R4KmYiT
e5ZJmkrQO6gtPlndGj+LCKk5Knfj9QE/yl0snuIOwXr4Z1Jg3NVPiXW+0/9NzzUlQpx7FnRnxvO4
STy7hK6ogSpHnMrQgMplHPuAz9Nv/JR0OIJmqMIiSZxQTGtKyOiqUUORSgWUYSQm98WOj4n31OtC
Edd0cEdA83MJWR7cHp5bAPO56/hZ/HRpT0mPH+sU+YYjCA3kzW9GnzwELX8irWDh4ee/SS/CUFm4
p/iQT2+/1JoZRyVKatD2DXQiZWszsyR7KzVPcWPFwlumIHAjM0exWOGTdDQcIalxg/Bkml/dBcWK
2fPaZCuxoIzTzkJ9V7QBhtfsE24j9dENMgjc2kZbbAn9wxh/zLPFWd734l5p6uxKMGu1kzEBjXi5
RlvRGppL56sfdRkq12sOJxryvv/NhMhqE7IRbcQKDb97OiKu0GCedJcjRr6ChquKTTOE5RQ3YEnb
spVPhrCMWr01+LF3DRbUK2FEs7XhS7Mq/E9C8vxds9xg0NWA5kj9wu+wn5hynUPchx4cgfpNq0/x
Ru1ioNGJ4S7E8/iwGU+b64yM6RlvphmDzIBGqBqz/gFOhxi8mCTa8IdeG7nwfoguLkcoVD1kum52
z4XYw9HpstSnGjBl140leBZ8LZaMNom5xb9omooeZXBzMRCBd4MmhEw5wEBzfPmuSWZbwlNq/6u0
Whr6bx3prBdjJ8IsYqutSPR5LQMTh5ap1dwTZgGk5rg79CWnL576J4ffY+RTNM43hnYhjTdwOTxm
nwvVeipgo4atu6EjTO9HxkDvpSdp1ht18LuKgP8GchSQOE//wzaecYJ7tQj1DLX8OiJlKufS/HLq
jZttJUAucUUfjjC4P2n9puJH1lKiYh0BuNafO0xV/om4wu2WmHw0Sh6zjsERPMJwomPVeWCmZ66v
BmgygtURxp1sKJQRF0bESTVPKdGTf1b97ZxJ0nrB7cUgHnE1KBWsJkJSOyqhtJgNOkU6rAPEAsq2
6VN64/gIc9dAgg49f4nUEkCfzLU1UpuJSD8A7hTxDKILlZftHoj69niCYSzdnvb5b13mltmDdr9J
uoLVfr1ioxJdfHCP15VLX14uTnzyWyVmnHJHc3s0tp6nQpeNj9f92RnvL/Sp+RRhPHg9/RzKLmq6
8EF6aGht0B5USd3EW2TyYpF+oExpLhEmQ568wbxy9W9ctDLuY57Q7VCV9Pxnj7rwXTnnlstM95yh
M+56MC+Hkh0qcl20BuqFv3aZ+euUcz4vIrImLvY06FZxBHWuyOe5JNqoyFsZMcLwn0vcHR9dLI6k
hnU/Ij0n0XS2wA3gH+3qsbyZXnMp+rOFwJ2m+Clya2iUdy4FRPNEi2W47rbLsJIQKK8BSecq9ixS
Sm3+MQVISU+lmOE2VpwxMgIBG3aETNeBfHCttHAt3AvhwMF9r91WaiKz9V6R9/OgP8ZQX/nYkLYM
tWFqZKAWZwY/56SCX+r0tIHZCAHcdI6k1I2AsD4hFTFJN9AZkgODSBCCWS7je0UXJDEOxXtfHKEJ
j+R67AWFu6Zk/z2QRF7w5g7avZaHWihFPehhGHkxGbJqRz6zUIx7Qx6f7pVEDKVy3mwbNB6kVt6t
lr49lhSCPE0VONerjCPsyHYgkFI8/Sg1h2D1AY8CgTIXLkmXAMk1kUEXVEtLslcd0TqyLm6mFLov
9MXLrSt7g2fJDRNByhv/uGTg62ioPWhbAwWhizWQSmH2nJVlZxkRgx9EuhGyxHmCDZQlApLOw4hs
dPqaQYVPpUiW33aslUIJgLmiF+ez4SsNtUAjIHbydveQSOSIb38lb0Owj40qy32ndMA0dciO0F+W
MzQLYoocAhCTZ6nQxRfooJ6redCb9GINm1SrP0+h2f+9qLrpjFC6PiIiyPVEp/NkiZt+QDLpng0T
9Hm7Eru1xIfMnK5iYxgLwtbqJTIfA8cgEth3GNYyDlJeAHb6q20TlRGBIHj8qiEpLeDez/qD9cmw
lDHDAlPQ4mRthDkUBVx5hYyHOkGfj9x1tJf5XcXAGYXRUqaDy4V61cUke6Jl5zTrZSRQ/mwyHKzQ
ZZybWzbIsjEfnJe1LSyYQ3ymRlyrbymmNiIBPv7W2NnbIUxcIIIsD3DKuC52qFtTgzXPzcpsRhL0
4pPuQY2TIc96OQgSizB5BmSpBXFSj3NPCsaEc1K0Enr8FgOgE8jgtsndWiEL0HxY3jsK81bLbKdW
MxfPya0aM8CB69zD364BuIzlAYQc34B4hxWoeXIg4jx7d0JRl4ZjTfmK9X4ykTeroJY2Ix7/mu58
38bdLJHMAHf+R3ETg9xz9X7tRAPskGVNwWxHb7pNwK3gnXEhGqVi9rhlod5Ny+5EY4wJzRVT64CC
9ai4yLnZMbOcRYOPgM8RWpricoSra8VUIsoGscIxjGbNxAAthaX+QtutL0UiW04kvejr//q8QoAN
F6dPcSKoc+HRQfNRKtyr3W1KAhtJ+IpQ7l/LcpGGsE+unt7C0/vuls4xdVntcOnKK3m1RdFlNo1N
taPFj4A9695EBO3okZvu59vf9p7gTFif7f+u315e10ZEYqoHuj/zdQ+V+6+RwgmmYr134e12Zw4h
VU2yhq8OV4dep37Y+KFt7CpER2y9Etg5/NTOEn5ZGRZZHiWIYKTQsbo8Wi81Zdk253uOCf93xdA9
NORky3ObvXINVokhsjq40KXEqyfne4+yktCMm9uyGbzRXl7NXAosH6vWQj1UTf6GuvPgqtsSCB1o
FJ4ptF3e3US3qvxrztM574Q0MK4JTIrjF4fIPTnBJoi9GcHtLKtGDVlMk+D/0FM4n14mANqRW7zS
QoL9V4CWVjyjiROmUqddFrJ0wLCa6mGyFV0OcQB++dfohxPei1I0PO2P+Y4DxrXTEeIl13WAM73p
l7snQWxWUmYLBYyZCxeSe+W9l7dbl/cC49vxQzpOd+WUuS88VIXVtI4wehlHdKlZdFT+Q9WyvcsI
Ip56ngYjDvxMvdiDqCi6L+eOKt1CBurFn4rEy4mtAtR3d+GPy1YnR6CYxsujwJEtW4+GdzKBGQN8
/tDP6VHy9ofWf8Q1A5jZ/Kjn7XrJA733NUibhtStZh9aBBMDhOpNFzzyH1v62/bd0xaGAHc+lwk9
uw/ruv71s9eckSArTYxypVL1Eeja7NvHwEsYvydNY0vcBf8ewUzRzwwIP+d6enD3l44dfARnSMI0
VyhEp3vtABcAOggAxW3cDq8p+hufZC1y5dN1GVDKSTr1kXhJ7S8O3u4ch64yxlQz73tB7ayQovNy
41sRXuaJ+bV3d56yJ2V2n8dbOVnWfqRh3MKg8UDsorYQ3PD9vfkreMegz6IRmtic0bi0Xnbwr2w9
qsoLxcdZDwyw7qrHNvou7lwXIBaonwDDcNPa5nNn39/P3PpLjMd42PwmAdwJaX7lQVhGBNLWK385
dcvhpAQQSfn/huwTi2beHBUobtdCc4OTr+DFEQo6r8UuLPoIERWtPOQzfB/ESKaD78/qYQBMQAXg
TRg1q8ZPQjc45Cs6vXqwisx0hGVSJjP+UwrlSc6naYNJcZrPovsW6kJYM/IemP5dHfqbCis3h/IM
p78QKvBgtUWKdbcIyeZHCbocBDp5cY2o/ho/fEo+b7u48qKwqBfc9MtGrs6oTkekJWnMmfbsvsj1
PRWcrFEsOXc2mgpNb6Q0EtiKTbCXxYOByaRNN7Zb1ghgxpexqA/IGYygZeBKpbdw1C++f1Tfm340
K8qDOXk0z7Wn2ID7i1xEPD0TrRfGPrgCyjVXs1k8dJ3Lppucr3jsZnLGOk5Aa2gAclUVczjrjMqS
BMmJrBcJAH4wCQkLisiyeE8ahE7tMRU+8nTC6z0bGkVu+gl8kM+OlYKFocBFCIixjiP8n7jbFkYs
57fTvRrPtElN20EqkoEr6GYxQcOOQtUbjEIsvvCDZwjdinm2JbOPhP501A+w0O4nZl/ecQiCb9wT
6vMgCMTJBtsyzrZfcnoSXkzENp1QoPqzCW0Tmp7B/TDmpz3TP1JWq0t4rrzSqW8jPU8bOx3b5aev
pzs/Ayt7pOUfLi3aZDtq4Hp/8xabFMetDio/raARv40sckPARCXESB4P2T6kTQRgAYLLO7zCkLgw
93RzS0FOi0KxBYC3YHmFy2GLCXwpyq0xeB+xlQLiwjX2z/4k6y4d5OqH6ITApqjWlkfTK4U7XcUM
mtKQ5hUwYxOpQGTYvLcSKAUaplfhAiTGPDB9NKbPNUCnbjsFnxLpMujm3BOOmjZAfJcgjjrfJD4x
HFP6jyeZKAIZCYMj9lvRvCdA5SKwWDIxtPhZe833cWKedWVWv0K/xWEtRvbvduNbbFcViXpAr9G2
+Bfqc8TKmJ5M/FFAVlimYTCs8oxxuHLenwsNPhtMVOCqYj3ZANdaVZqWcStNpd7hoyRh0kxrugXp
u+wX+ZNZi8M+f5IqZKXHRz6FPox5PPnsIJR0kUSwyw67acEQM5HjveFcWi1XGdtsq+ZTYESojDAw
A0rkYBu1hmS//QFBHoSJkPWqywH3/I8frV3A7LjH6wKO4kYz66iRFelAD+DFuxcAokktFvyhgbBb
hrSoFvyXg+CHh+4yeh/++oBIv2PbFud16DzNhrL6kDw01MtBt8VdUknQUlrhiY6lxgUM8JwXH5bb
f0AQYw8ou/oFAE/oFMOlq0A6wpJvmOtlkEyFBLvsrVJzs5SawQfSlbLj1Ka70wWwZXFU9PhEP36G
a8MP4Sp6sZFHlARo2L3/y3XVR/nHJk4aZssoiR5V7u0BBzVKuELO1kmWDX/2KCHdsJF12+OmqvNg
sFBaiS9/L183VEm0NYniD9DUuQ5hn/UQRm0ZB0HFas8P7MRaYm8d4AnMxMqY/xVQ2pkk6hNeOWbZ
oEbXNEoXEJ1fUHx9rzVJQb1Uy7f85/IM1BAhG0P7Lx16Yt9NKnViS0BP53h7GzVwT3IDJBAvQvBJ
Tgr47JrXW1An8wF9mSue0puZH54Rn29DL5+eXGr7aPXNNL9ud2IiWmmPZwIdFiA9S2Hl1YANM0nu
y9p1FqKpSaLn9eH752CbmBjjnBkeOpI/HZb5ITbjLrntmPXffes7lAmlwfwHOeJu++L/hsLiI+Gi
MBN6njdQn9IaYwOidaorOJj92pQDI6Tlq2kuNnQD3btBMH6odFcULd0hom2bCPxrUFDdAWmtcOhV
sS7yDOrWg67TVTSRpUwlzktxJqWjjPPhK1oZZdSgaaELdG5ALi8bdVFzBVQDKyMd65QmKKw0I81A
AWV9B3GUeP2CCOC3DjpgCSpB4H7PPr47cqwhVbuoZQGf5M/gdlmFFEGKeFwfdn4Ib6k1vRBxLNwm
anwlXDrn7wBFQfYdJuKqFWmrA3mMYwmBrHenN6uMbSJZ5gICrqbgWAfDrTcZJyBpJ4uVyVYpT96I
dgQc17TneEWqx3i6nJE7uzAT3ORxWK4N93SN9l6hQK0eWhLqfnqRK/WVy7X4RC4eAzQPwSqhiq9c
Nd2lx/ra1Je+ZaO4U12mS6MkOeXA86XnB3Jh2UEZjdGUiKtzojj3LXrAvCgnDMkviSTJVjUipgWx
grffwNGL6VNFqI35Gnw4AZOVyUgc+gEoeFs6NZMbunvm3B3ky3pHsoLBPTshu8dVSzT9FrzFv8F/
nsGeokh3XKPxqbD8jkPQfQFKOWp8pnvZDAdt8v9Pg9D0ZA0Vg93gPMEpuaWomf8l2oGY0j5UU0+Z
dX5fk3amOYDwjZdWMoWhEESoex1X3zZKu195TxDbtfCqcx2QebDq9N2HlCHB/90nvs0uOEZMpgIs
1au/3OS0mJRnlf5CFTw90xtoq0OUvzNO/361hFL2loKezOwKrpFfWUgK7TWpi5Rnz6TzhksHiqXc
ppCGFBqIe1Siksg28fdlpFcPp2x6W72nM3LVEofopDageLWrUH3kfvNSdv0v0SUnTOd3cc6SjBuL
24aMSKjkRbfZz5XGYg83L4CopSlDxwXOk3icerB3BJPc/GteplpQsPk41OkrmtZCatMF+T1DHiGF
wGBIcNCSv59NoqhD8JqG9AibVT+9fe5LSsOVOuPJVeHgvZVYQwdAmzAi0PZCG8vI4f+eaw6rUNYl
N5cmdZkmI5HU509nXHVvHUdka/NU36Mkhi77n+YmyGvYS5eAT1PrLZKY1NXzPN7VFU79KkR+2h0W
rJoAZWKdCywyGIabw8ax6tnA0oY3TWuFIoQIKat8Uzyv/1L99HQQoOQVQ0RctDvDpSOclSiBc4SX
+kFbLzYzMYil8cf/BoSW6d8w55Qv346uAb4FcdxK0z9d8Wt2/KWSYt0NE5quPEx3jWAy28NJheWW
PqY1pTihILP96/8IR8Kfdf98r8CYCu9JHjiaIFEc53vL5tVz/8WdVyLifMydaLg7WlhTQiaAj0kQ
XaLd4peppD6NpP0V3hfeuppcGbrA1swjMg4SyzDM+wcpQkqaVKTPLeYp4XScOoa6OxVCfO7ybuI/
4gtfIeJzrzp+mr6/PAvLlglvF4BbAyWdSkK9w2JE42xDQdchjBT/GQeWXVlnC+pGpeuhhAwiZmoI
eYJb0e0wsWU0y7Ramk7GZte22qZoGyZe4B6F6uwNSLqexxylxtMNffSuB6WUkS8aRrWC/KXSWf8K
huiwahwZizuXRP2tj1an2XDPF8V8ZQp92UQxn25ZXfyrW7FjV2A7CQ84S/8o61RTk/IRIPAZo4Io
i3ZTEpPLY3vfDwEj2XoI4lk2BxkWO/fWU2aq+sPbyqaWwvsL8XZn+4Ld1Oggi9J+Z3ianUG+lOtJ
WPIt3CU4YyzzqXI979iVyObFVOkKpfdoG9h7A7ElHATAMnYEydk+3Lj7it1WkxrODSo5dfB8vNzR
yjznJoMF3lGSY3mw2P9gHYcWD7to1hIAIFLM83p+oOVWYEZjh3gHS0EEugIBSHven92h1Z/dTjwf
GV1kttWQWBglqKLrJ3LrmdhNfn6BbakzJYoiKhleGkEG8IcFIadlbujHf7NSQ3gCFTNBJy2ElU/B
H5rmMQfpy9PywBEudV9WSzvfif168IQLmPwsNen9Vqw9m4hpwAHpSSRS4fE5nBKmvb2jr1skcPc7
PZKwKXrH7JKXQymB6B0/2RwYIjKiwGTpQUuD3/gcgA4Ymrw8Wihks8LJvOdNwWwx4AOy1WWSvZ5O
v03Beo6kOIINA/YmGLCAb/XiLuO/PkLz2dMUmsWb3es+CMuU6Y1qnZ1hAYdSzZ+9jxhJxJiUFuc7
Tga9FeLU/wFP4mS4MCVH+Whx8Qjmr2dxJWFSd7lDG8lE7Q7MhsgsUVRubrTztIdG5aAHD3XbvH5K
TUQnbgB+uLaBVHcmpy7SCm2oyRx9A5vjvl0+QUxSXttsQE2Jr+IedVrcCiGd60xsdt4QC6XBqu/4
oMIEKRBf9Yt96+QRbvcAs/7wfY+KbHnRGVjNppxLR4R8Mf7qPYW5HlpRKAWKms7+G3aLgMtS0pCn
z5JeVUib9d/1vvs7ep263TneqhAtn8iQiwsUtE9OyVTXmhIZhacqAf0DSdesc8rDlem0U4r6nOTW
alGEtjxfGlRD6pJpp12aNcca5O1VQH3NI/ztMrzAPavY0+BX1vqGPFti6dKYxXkckRnfzQks1x+H
x6lUCxbHD+PAd8ki28bVMTSro72BO/EgF/pfSAkBXy31tM4obeCkOAl4bULV8Jl+kBVk3wEQj9xx
feEmogGmyR6YSR6+BtZYK+kC00igzYH1OmZlThDfELFX9qGhr0ILBohA/MlGC5Eo65fsD4k9Fu81
5BTkhPkB/Rg+FSqp+ClEGEMkfkdKWnKRZk11MeUeQPt4VNHJcWzr9d1JNzosJg/eqq5pc4cGofcQ
fByuTmEVEbMEmHlyflKqmhxcENCGSlu7Gm0uGqluJhAcQt0IU/p6WxHLaYHEyPhToV0M9HQqhSgR
qp4TOOFUAIelXjoARO9Em/tztuYlsIns7UUj4ElyP9kGU8VXzodcBGe1kMIG7IGhlgGo0j5Urqk8
NwMbg6ZD9lW65hD9d5bxm8ovyUSi2Ez7XTYL2fLVAG9XyLYEqO56M1wpnih1+LOPitSunWZ/3NhP
0y9nqjYpT3AIdhSUc+0rE2MR9/3olXPp5VRrz78brCULQ+wpB0fDajHS11lA2tymwcPGxoBoZhda
DMzY4Ane0qLDkejkT4dOox0HKU+l7gKORGSeGr4RqhRmrFCpdP+7jpcJ8baWOxzSYWRyVROMtTM3
yuy5psUYPy+1pnA6uEV+4r2F++Ls1+AzOd2qFcIksRdW4LQ4LHwKroPK4n9u/xrLp9k5uMmf5AZg
aMjSwduIpt2U+0Utgkt63jDPDiLgh6Npu2XCyEFm9y43WJ+M1XGokajF6F167Znc8o1IPmASbaaz
PlwdASIFM9G5X2tj6G7ADViDNEFhjwal0G0ggjqc6qAyDXvu0yBIikGSZ032uN+ROGUIFMwNcCmm
zTA6r1xvOYWka6zx2QZPIyFOD55V3TSCixDl7nk2+FG9Nz5nrZyznQqvYwYxsue8Z3D/VDrl3nD2
Ncc5VFVBJXTJ3LOR9LRS+fKG51CyRBdqfR4u6DHMvV5RcbA/EecCyCM/pgiWARkY+ea5rbxBE+ta
G5B5kMhGvlUdfGSn+qI8xK7bFKP+qPkws6f5JcLkJNdO/0kD43SLK8Gfxf89SmGWrO2oJW6F7i/f
RZ8y9hdkqyiJtm8Z0OcYtgqLmEc0TNZandlj+4khYTtW5+2GPnHcKILGWJZMnUIQNFhGMqPd/9NO
iq2if7l68WDOmRW5nJqhp70EnuFrb7UiP0Kyu5aDSha6P9qyWLeoisxCugyUFUGgRcOy5KMn57z7
YkH6Q7FCYuaKyslxAV1esAwghDUSI+PknD/HwDSJqfGIuxo6vCADtypF182EihElxVkZFqdozpuS
00KEh84faNQUVUgifyGCmD/UUs4Mt1K7jfsq3FRfg5EtfA4P9JoVbKaVmqOmjLuEcdgjOE/jQtib
Ryrh0hfrUdwdx3tnkY9w5sjTZhAuoQi27ijilIs+VCryJM9Be3A7eYIJTYVqT5bQaksW2jqiZytb
oeAqzj2Ls2K07MHhSFkd3K0bm9rYSZ9D1sNpxi7b+LG/Z4xAvwtykezOR1LeDZJn4qgDsfX9wBC0
LTaAhMF9SfiM6X9VwYgzR0AYOj7cMdLQ776EnDx538NMiVkKYNxe+d+Ln3mKPYDiV0t1pQ6u+0NW
d9XvMqy2YHcD8XJtQLsJeviUW3G9XvzsRZwHllA9omGJVWNJxG20V/tJeBWGwu56QE7z7Uw+eq2L
3tr4XCFBjcUR1JpcjXqBn3Ryq/8hoAJ3geLofbYNjNrlIsvfcBtPBoiiCNDFQpdxIm1MJ69MOdgj
io0q+WME4guKhcJpmsG/3BFxIPY+8RgAIZk7M0FZAgrA5PYREIHitCd8b/ZSmkrbocdX8DJIgbkE
fVF+uuxNxjMafTxJ9sDdBS2r9mBU0F3jl9GL55HJDQCWcveRClSzbwHVnwYxJGbI+iSrc/FzTKLd
3XivrK788m94x6QW5WOZV5O2nyvM2jT5bHiJmHvz+FSw/yU2K6ifVxMJwR1U8iRXrcn8G5sv5RnQ
rdiKI3NYF4uUIarHLzpkMfCDez3HS+P3HyFNR54Riqkdyu0M/kUn5ozZ0rE2s1JsnxCTOPEFaGEZ
zt21bv3LzS0pnhg5NnnYxhhYOx+ccxqNxiQtyihytTYuBnPvsdVui1/6R8tFdiQqn/M48N3TfAr1
qanJoyrUOCUVg5Zd9UYyN8YGeaYN5tUiH7fJ8KanOwSp5c0FPyL//pvi3nxdono1cuVK0W/zk9+T
0OXxcT6noX/TAdLyjoJAbBbJUXrTplX8Vh7sUU4REz4rY+XeDpyjoPZPF11JeM4B7fqjZIc9Utm5
E5bLYzxqkPj32zcsl+92B36EwcazTzLQ/SDy7sqykxqghOdzTQ5U0sbW7lB/pMIr7Edbrz+moNxq
PVS5/cJhiMaV48+mlUx13jbz9ozVTlk7110yvu2Ts4TeYWHc94luFvYMKQMYsh7s179uisvk7diM
wAwY+Ka29dOI1IOm/20HCkGPmgDiHzqO1g+3MAaRh9TNpCHXXU35m3SOGL3X1psJfj1zRq/kxfaG
ajy0CSL39+cQvg9OY+xFdx+1/nGqfbNUDoFEGR6/lPDAnC0I13t5V8oARHo9iIrKYruN5T7d+VgJ
10/FLjW26t4FmCU+g+Eeox+gHBUuDr6YB8doM6dvsDvrKGtIDgEhdJcqBBaymP66mmsr8Eczjz3q
toDaGBIYS9dK0GeIWdK0tXEAsePERjCdapbnaOZ3RLOetAfkLLXuy14dtw6WzdEX3z15G+8ae11E
OjFbDy0HWTNByzOfv7iGwP6B1fJW7pwOdcgD9UUf9S8iybqERyWE74xBORQPnmOmMY9x0mhJQFbG
fAZE2Js9sDam/ZICbG7TNqdGlCGoL43Sa9ynRvwIswJ4SPysE0F+f78s+cs6jZGA2EsLwT2rm+Di
oZqkUKRpREj6j+tCVkfLEyi7An5wwRIht44wp/OlU9kkhZFjadUO/0URR8yWD8Q6gQoXzZsc159m
95699mjwsfhPAzAXfXgBZf0PojBUTtiFV3LEtEdAuQLHZ0iT/QzJseGU6qlfZMgGZ7dWrlUg55U5
3cZtLs/5vpjj7MCQrDQKLQPwz6K6euI1ZKzfpLtgnJzjHIBHnYbnrAWaNJiY6P4Hg9wzzzdmdz+2
QOolSuMiI8WSec6+snPB+fsm2y9YYqPPOGltmeTpRIenpqyZ3Lm/Lkk8oveaIujeMrsfeqbGLtCa
hB7bTmBMBIWMjbQEDv3JYUf/BeX8pSb7ulpdabiwy1xvkLJJXt+P9fGk0+LM78ZcM3pG8Yj9Ir5x
AU4CiXvVcFrU/pP0a+0sGi7LW2h11P9tgAoxdDnWn3TfWNvkOvnMedszOQvfPT+J0mSFjGMuSgb+
VkmK6qOXubpVqUSFTCdMraRguaAv/GExfKNuyLDO7rj2QAsCLAWh5nVkmh20WFUzYVhJn+MElQH3
3o+NbZCNOIyIHnC4mu/OPmFF7VOtPyUQfRRxHZFaACiDKfG3+Ow97Jcz1QtyIspx6MNMmEXnlks8
38F5bN7CaNFd+3WWQynHNo5com9u5CdV9m4xViKapgDM/Q5YSolGRxWbjRBlE1Yx/2ITdF9f8r6K
pWABzvmcJlLaiKpZH25ugLIjZyufZi8wAqdCPno/HgZXTTYDkmmeEVtBGf20E4duYmWLe+9N7mmK
ixLGE2fNjybP10cfwIKuUtaVnD9eCVgX2kdlx4OI446bKeAKhxrEEIwwJL7eZTQ6WVAlEZxkuSKJ
twgKxzVYTkgN15HF99hZxoiOupqAJbm2L2OnEot/S2o9U7cndKAyiBqL47wju0xMfm8cRdtooysT
dohelPBsexWGYoQrBaSz/MDQIhvXae+zUuysE6jjFTD1UCm3IlZLA2Kh/JPD8iMdIjpPjwmaP5Hg
VHuPWI6U7x9D/IaCSzPhGAo+xEuJdV0PYiKUfFRKrQJnkG9zu4zKc8V4zO7qwPCxRe0nUUZjDQ4J
nKmWVQOctv31Xws7U2ex88Mr/cXc/+U7uhc3q9WrAuddmhFb77wx4vxRCbT1utJ+VCG/oNJVyfg1
B0rOXjd/wUM2Ru0z39ny9G94Cz8D/gwKuaTV+aV9RDVK7BGtdcHwPwK05aWPYZ8ll7ue1wCNulAl
hKi3Q8X1TWrjYiMvNRsmdqWpdLkS+gJ/srdh5kqvhJD0CFQiptgzEjxZ1GacdDOkxI+P9v4PKzMw
KYBt2HbKsbdIwGwTwyer9xdI8eXaOnf8g9oxTI/AmbhjAbjx/jRV0mB3jrLEcR3P/PHpBwAzxpDT
9DShHNM1pQ+ThaICNSihthHEUKMfmm/E4kymNQsJX0KYjC534mt15d3Z2dIxsnMlSjUsjhHNwtI7
scM5jY2xTlwAHltbl3myGbfc6xSJ1ggnkNxG8UuRRLQcrBkqwsnbC+VRBbrTbZej27TpHF7yGdJr
5I/qAkorwgtVd6Xk/h1+dU4rxn3WUHX4WotL+uqD4y7fN3rZwXcoN54B92N8ZioO5jiruhEgg/WT
FSMHWScnRIFRKus8hHhmelIiMWWaoGgZgSJjOjKkkVkjLrAGw2vnHf4FjQVmXvWhzm06OOuJO+5u
pHqZT7LpJyVn1NaFEtd6Yhj2nYs3mryCE7JRXFU7OTAk47CTz32tlzIUNdIidgDBcu+kDh9KhF1P
eVvNUvnOpcaw1yjU5a+Bpf+Z5bjrGAa3Ja9xzPIVlmtqtjdPKeUB3NSZamkdxQots9G+WhMP4Qnv
gMDjJhq7l5Pzat977+5IJgYlcA3OYXrWJ0s552xu/U7r13wBG6zg/gkvHb7Y5EiPrmT/EYY/5MSc
mYY+P7B7IzwVe2XxBfaJeK/6okfO4MFPZFhfU/dIqRLNJd5kk7ICLitK+aO6WuVyc34l/0ElEaJy
b4EmEi6xQ/I5VhfaiBIUkfk2DwjfPcshAG0k0GEFTywu22lLoxFkgpkg6rBdCgcnAueDsb55JGw8
ToO1HMZqPsnsY0oRLXOr1YVHpRa1Ci0GAeY8WyRdg/2pQ0doPgq21KxM8YUwkc3VEbqrUUNNZDnp
a9TwcBZN4UE+nj1aZKSDpyuh/Ho5j/sosVplkBBL1iQDrBZuY6uNG3miCNWN/uu7V6e5QxC7ryc9
0G7Ja1BKlILzWywze4EzrXFjJ7a3GaFY3a15fYIVjVcuFpAxt4ZIqOk73usOTb6yn/sitU1NokuG
2b8e1u4TqjofUChrp562YdOP4ocGU1jCN4ipHR005lAFnO/RVJ0TE8z3v4s96T/SnznpRrDifJpB
o2FkTc5aE4TxYMMcynt6zNWCOudmYZgvOlSf36scT7FfbfWWLhkkP792gOSX++yGdP1fqvY+G0/q
nftQ0Zdr7TLowHI5LyGQmNlQjvwSqe4sJKAPpyh50U2/0jcA34+15lsSMh6PDhRu1411tqv/CFjt
ERYvuUnjTWQoCu4d7fueY42STau+TLo2U2C0rt/9w24QlOzMcNPiqS1iOVE65LvIYEF1LCScRN8r
Ti+S7bUoPeKY4OPoQOUoTPJAx1E0udvPJ9QRUDo8Nq4+NnQbL2v/eZ/znvu/F99swXDbXFcQ9BIu
LrRLpBjtE+LbU5Ikk3225HUDThFThhpNebYDJbGpg3fQuiPwMyUHL+ro9T/mKv35NR+KLUuljd4L
5BEbKDJbjJHCkGZbpoCk/IT51JCj64hYJCii5sPvLad+QgMdeUjptVFB9I4+bQH9K4HZGgHTH/Ru
Wf0sUYlq5J7kPlQfcaWHA6LwnicWKi0MOBAWxYQD/rBUDVOIVG2lisfl+oW8H6dxb5ULxk8NJdfm
HcfV7Nf6r+xCTDBpOl6m8hzIBeslNtyOhFYy05CBFVFzvkGYUBofYjUCNSnnVN0l6hdi59ROPFTH
d/+3XqDlaQzpvzvZ/VVpriNQypgettMVyJs273Q/6gzPChFMpC5SeDER3U1RKUmkPmiZLshl78/q
ht0t3feimKNbPKVjVlUSQ2AQuimJu6rFt1N5dWt4p8bupr5W9PcC2Sjzc+3BMW2VGWI5BdNQtw14
GjrslejKXQzDoc5SUSd7GcwHvptkBf4sBTwUdHcuzKzO1xQCcMNusSma/UNQTGwlL8jCz4mmdFQs
3djfdlHGfItyqSmoFJIJanUzRwyL8usN1vlStPz71svTdpGMl98EeyHOMX4z82BTv8l95tNIV1JY
LNrL2eQP0MvXW/KnAhTtAxHRGvuQj2Fs2+bGflHch2yfbv93Dqk4BKh6ZTBJSRoJmRGc8QL5wdCL
LVD/iNS/Y3cpd/YArTV6CH7uDxHwCeGB5o2947cY7VGA4u7s6g1cbTOxk0aoKew9riTchut5SK6V
z4zanWlh3oE7HNs7cErayh+e3Y8Pf0NsSGxPyU9bSsqmMZmBEIHfbf3Q2Cncn39eoewJlpmXGwjI
zI9sD5ZDDlcBGfYNHL9XoPSLs2NLVF1Qzpa94g9aMEO6b29ujnFLF7eNaWmjqt25j74kFRMk/NaO
aUkow8MIViXeLfvFe45k33RW80cV/hp1LB4alNLURCkMeHfxGGaJE4N83HrBEJ442dEZ+1clRMs2
tLUsFRrpHt5o/mnlDbr3+J/pQTT0v+yZmeKzU2GZ+0O43Nn4nFv7GL0ThLrMbkDqRY6LWmyXNjxD
qoGyRFrXx+2267iosrslgbH0R5/iq8b60BODnwkOL8tOqMQdA5161Aers0GcR1fgSy9ey4ywqbdv
d6vweE6PlT17PiJi9+boNINlW4kPPRUFMC6LMSNffon/NhzonunN8x938BM5nAYErmduhzFIdFKa
Yax+BPsVBwnYZiyGifx3D1X+CvkYELfKNQ5ALIKlg9GMTR6L1NeKlVGsBlgZHGr8cVIes9R3/Ai6
XBt4oyWd3Bwh9xnHdIXk3N1VAL3HPxXB6uhjXRpg9QW6FogMeyjBtL5KDvKG8hg/4ARAsVw+1Qv/
9rW1TYeb7dO640hAeJ0eL8fwbuymh1iSIQBccWoBdghW9g9lr0l0HS02hcbvbadSqwxi8+LPMX5r
2ok6QZI7pnVq0GHwZBtPTuHm3ygP6fqD4xNqB+mPQ7LNfcTt3VCve3FMF1MOQqhAeU5ubfJ9M8tQ
mK1nRQgKQONjBDFcV0vQGpRRx8ZLCv856DoeiYSAG+NkCfP+EpgbTRrJVF7q/y9S+cw751lrukcV
DvkkvmPVU0ICP3NEUiJAoPstJu7qS8rqGkDXZviNGn105MlK+96S/VjTGbaakfs/nEOKFBULgykU
2cMXIyQ2+fxBYA3vC+jjA6odtKscbg7yD8y04Zg+KK9zBe54edvs4Q7ZmKlDeVJJLZ0AGjg0L6dl
xJ47avH3y0GD2GDoC4B/RFMElId/C3mWi/EZiR/T/Qr5rVazIrtuYkTkihXsCOrP6aaUgeaU86Sl
XU2Yp2YKQ6jFP+qKIliazUURRzJw8wL1ONb8mY9w3gdUZLCsB3sDjkw4bGYxa8m0lMUg3uBAMm/Z
szTMUVOPqYyzIwVV5q8V74kAsHfCbpeVF06HJ3MRDVY5sPIFnJorkLjUsbh6pXK9WA8tYIs2dUrt
sqyQ30Pmg0MpA8wmq7do4aeYDjWTZesVgrJJXdx5XNUro0/2TelL33eDHsjC78g1keopscNxY1Rs
Un5gFDe50YApiLuI5CyVkFmuQSvlwpKjMFV5MPDfphfna9YsI7N6O1NNo+g+yfrHHVnXsa/4BX2+
ixImHl/q432oQwWMA7oqhAck+oCZyj4lFjYDRyt/rs2SKvM+pfFBYaSoAMH5AHT+WLjJWAco7R6E
HX1T7Yywf6tphkW8z6NN45PC6tUzVEsxaUCkq+57ca3xJHJzEXHY0QPakBVdZkI4depDYqPHNNxr
veyznO/faWKqUPawBpk0XpLTqxPkwHfeiNurEL9SWfQs9ik7yu9GbElwNKdBUkfcVe8sSSW2jxro
9hcIqm56wgvM4YVQnxqwPQWqKE+g1571UX1RXOrgEa33GOArcTf3J3hMnpyKy8ZHmO74n63Be8uY
T56tX9AYjVGHvMZ2MA1xvuzYYldzUdZctTxTyIyCJHoih69ChvacGDNWrusRqADMfoAwMloqerXE
a6TARxNo8dRjgtrRKMWB9aRPXpDxogZSElIpXRUrY9UdECT5k0v43XCjK8uWaEINTH7UqwBjgijw
83h5jSXPIjWY04MSuNhurLYgMHEZ/ry0PNtJI2EXFLjJ14IExPboGyIrJ0U0h8tLtY0LYUFTi4Yn
c+US8C6bRnumG6PpDhLCQLyZSWP0wFGUwT5ZZyvDI8NNoG5iOa87rgd5gHiwVjWo19M7RFqm/tES
7+/vmrWMB/eX6UtN2Ws+oEtsjPL/j3TcXFF9g0nuOr5ywNm3joEWHche0pKw4KXeIEvibTCxHlGJ
zGb9ngl1QAGAPAgVnT9Su/eULF6IfPSUde5rLHKF5Xxy8ohQSkP6b3B+s+96a1rBeteQaNdeZLsM
phRXGQMFEGICLjfkY9CF+UW8/VsoV2VseYkr1SNdrNBAGDvTWRBhGWi6bBkihw2735GPaVIvnrhT
xPKrNrOR1MKlQoVwgq1GcnEHD7W19/SlvPDIVbh2FHDi2m13EOOeAVCz7bYZi13WUrtWB6K8Wy0Y
GR2fDXPTPkocmCrdrxrzc9TuLDQeSMLuNR+DvFngruVAssNPXAmxy5WY9ndbpovcmaeUNpXnuJ5x
pUmIJSPTCaIaNjKC6ZJzH2/YG73PML7km95n3Yn5fqZ6A9Zizpt5Cp6vy/6zcFS3/U+ZWAZjzK01
R08lfCYtcugVxAPmz66iGtTPX4ARWLVW4nUmZkaa7pl0tgRzbPNPtjnl9UYgmg3XmARnF2lvemuI
ifnqZAqC4xF2mUMAesg8kwSaIlEWJG6DKFz+RWmR+Qxu8gxtgwHuabnWDKIhLiOwfqVlO2jqfjrZ
5s5wSIlUz31iTqnxC+YgYM10mYhqk29d6BW7B7WLy8KC5JAMntIF3UlHkDgVQl/bMBD7YSiVg1aZ
zTWAR3Q52hOTY1tQM//4F6AGptvYccbVYjlvcBQhHFgken80S+i6yoqDVu4FPf6IntfE5hx7gu6v
TUbYk0TUNsau+ADHLp1bQU+uH7S4Dw+AmXgftNI61K4k5ruXQPWgWzka53XXu/SqCxrHHOZY7uws
AbCbLFT5s5KT2AxghnISlp6/9d/GcDkr38avHKEpRCiPE8CwLT1rvQW7w9tH46qCODshAbuF9Pp2
Ap75emZrnAdzvMoD9sXiY0gcl1wLumX5RcxMMqHqMw0zOM/ysdfevI0MLBq/DmoNt2yFMn/Kggwq
Pc9wYvcRW6/vtLwPwYk/0+qeIz83auErbGmIpM6PzN2PiKjIvSXdl4tGrDjGD/ZABWTM9aKuU9m7
bJx58fK4BAugtiHZQj21LIC7bO19ZGipX8tqe4XJ55lGgJ5gDaSBYvYCDWuD4us+mIgzsb5OWpk7
SjNoumGrSFfy07u2LfrvvZogDLB7dgt7DI4OYvJ9yisRwZWqcrCwajuPeFp2h2mD8QG8cYUHyrjz
iNrgnt/WDRoJOAyMlARQqU8K7D7qwpOoMjhyjzFo7NS0wqc0sc8hRaHFlWxVlVzGQjT13L7SJ9lu
rJCiGxD7wQF1Jy8+69knKH7oYtRUdLaPW8IcILBF0zIL63pIHoVdunT9721Z08WVA+WvCT9KjDAh
qILGroltgYgR4lrj/oC/c55FmRdfycCu6J+AmE+XdMrGrzvP0H/J3duZQhARpgphBYsaMf5sD82m
b7upplLEP07hpBphA7CKLJ7IKxmGer/dbI2bZRyM+SDVqx0NHwdF6eO95kBdXqf3ucggxTvyEUva
eCFE60Akth45R3sXGK0JvBMFnFEckEZ1fXFTvlslevNoCLbQJbsaRzCfODI2mFYeOe1AjWExguyM
UIFYBCFZ49g1XCg3ZEGNHHOJEp6gjcanlNuf1h/1cQcm6qDYu0ollj+JqpXmG5SLOCr5QqTRHgSJ
cK+3I2RrQaFzBIm5xkfKVpStZ3tLu4GyY816hOiDEdbh0V9+1xM0AAjUvzxw6V58NfBxD6QWIY2M
WVuSNZM2Y5Y8JyaLjCYdililmfNeHnvM/IguGs7g+6xulJZDQqaJ5mC13SmnB+iTQSy6vX8ryjf5
TrQX+H+/BLa1DQx3fAWhnPkr31j81icTZ0so4xb9qGVJfE7JtrktY8XBtjulEMJJLfP0/+JF+sM1
8wXu9Vu26Tpw/99EJzR1JJFKc4bLk00zV0FvDhEXI8qNnU1v7nct5puR0JDct7rWX/vTuY7DB3GI
+yZwsKggVhoudh8Iif9tapCCcdEqLrYAYk8qbzHYhCKtf8TEEyH0PK+ffP79eVM0T4n2u6F8qeEt
obOSawfvv40wJnlZq4rA9kMFUBQk7n9KCHiJxClGSlsdDJgRbYyvqFeLXLERCxIH81jCJKCS7mkA
/wF4cHRkgvhl901XjHSa5il0Au6nUgOzA6HM+cQ6K8SEG0fLjdJa+Qf4/jPN46UaLEcc0cFba2F3
oscYdO8v1yEigVr0t9EzzFx5FV3ZS/AV0DeWgMQGGWfR6azOh5ROiSYJ6yD1zEtg3qhCWloMBqss
+1jrRb9pIuJzJTwcfoioYIPwAXXde4pozr7M1jHhdrTHCvBNyFWHImMaaXavrvZmXtAy9r8Rgv0+
xjtNAQ4BWurqU9AjP978mdFl3wFolPFuwdHZGnxPhA0YKlvsJLeGq65j4rzZFiNN4esXsQ2pfoAr
v1TJ6UU88A0Vb8yXHeoCebu0Ha9JnqC4wGTIwSt0M2vXVIfvy+z3v/QNnxIg9QQplN7UHhvlllkz
ztP8HN10iMt+WTGiUYh3I6jRWUpEuOPWz23KRH6DPkmp5jdG1Szfv0zAUy5PiQtSldHcEbC1iXSv
l//EsMFNcyC12t9g4egh/5iBrsj4zeXpG8ys3SPUxabTAdB2TpcvVbQmI+8Was/hTyahVOuQn1HQ
P4eHhFka3nAK8KbZWagL8aN00WmbPHSKBYKyF7hjyGHqSwalXFnJ/BAepwARuwfzRbnE4dOme2VU
JKUqhztDJyCl+fFijDC1ptB+v/O23xLBdEVm7xWp4xnKrN3RlnsdTQ/tQtQ6/2kVS9M+P8M4R4kp
zRNNCjslweBjOOh8Tp1aaZ2bK/gVvZuyF7wtOPUNxdPEtbV6quZmC+6XuXcVdLbAiHqXhCqMl45m
9+JzS0PwCufJ9sKqOwbv1cdczK5SbCaPmKH1/7cqXBMQZ8mT1A1aXGSo2Imvr+X6l9FyimsbMdsX
OJWG51wMJUE+tT/8HJwEWTy1s6hD/QcP3SbyY9L8uf5eRD4SbpWKY2S3p7NyGfGsUiUPGBrcurnP
TesnByDlmVk+0PqhCtpTtNYE//NKqvfDSfVYP+SrN5WDYiBWHjOR7TS1MXN+4kKFnOC8RJhgyELO
VpVnWS1idGT8xJ0Y2h7Wd9Eaek5csurgANCrUhXqx66giqUOPHBNbdbuTgIeDd0sKcSNDigXGWQA
HXQLzqSBBLvkzZPg2ifOBoWAEuvVxfbL+TFgvvnFfG0G8qpaz7BZlcE/a+/poF4OVSVtnUEe3HJK
4av9ttWoHG+fz42QpFgmFJhRfkdTX06hx7/6R+cNqBxNZGq3iUFxmhZesrqM/pObCRZckY+yiC/R
3AkoEfiSHhosPLzwCbcvilD4wigTTJc+RQ8xZzwM7NucAmhgY7vCueCD1xh+iXV2z/MhR71itMj7
EOnZNZmOr2fMJZ/gVk+Q79HRdTcUr9ZekiETpK4ssDuj7gmQ85jE5UwEuRv30oaud83D4F386Nzz
FKSu+2JprDGPwEewkAjPehpB0ODDET6VsyU5eV+RQIQn+Cphf4vu+pn3RQfvq2kvA4P5S5//onXD
6Dkrm1H7sIXBznmF0Y44UC597O4D1ragnRSuWx8TYfMJTxopZzXHaesGQmOi0LSq3w2YotFuOJZ/
TroZDYUaleJwfpAAxCBFaA/QDul6bYGwjv2ZUXZE7f5UF9hqvTO08Iqt69TlNBudBe5dxiYyT6ki
aXIcM2og7/5XTJbK107iWXWo7xh5xTYJWukT6EJYV6ZIFFPoHUH+32Qa1pdkFath869tgA0AKPHG
J/Odg6bBK7q82eUyDzsE8eaN+j8iA5Tg5P4PA99Ixo0EKe3/UciGqiEaxDtzuZ/bUGl1DZZ2/NWW
ajGWSPXXuVLFmOI6W+nVu9Xa7uen7CU3w2nmPp4S8oQtLhVo2ZVvFE/m9yu0GA1sMjf7G70EFwdt
Fx9Aq5X9uRdVCvvv+PEVRQfUTaY+bRB3YunfIFndso0lNyh1+O49J1LbLpAK2ucPRd8otodtbwuK
LLyMVYlR0ofWOrm9lSXD4Rl5I4Q9Z4tp97SFjD/l2ORR5rcbGsGUR4kGKOu39K9CLkCqod+vQ6Yb
abcHPzkTUrL0DeUNBHTMbJcHSFv6P0g+gbdm2u4f6cJNpUscF1mYO3bl/rR6MFt1lMONURlXtC89
oBK8R/OBpnFTZ8h4UtwSUR1qSaXWK7QOm5AbZ9oFxObjBzWSqVgmpBOzuUcqGWiQoohtofDBXAiu
Hjb1BsXm/pLtir/QIBaAcCDje5qJMYYdvxI7ULoc/jiqdRARGbZFwngj/CBtsZ6Cvgb1oMZJxUNE
iLPWUslihbz0ch3eyez2wMrbDr3MHJ/MguF7zJR8bRmDQWq1/C9ZsLBGV667ztqQD2WydtJNaAXr
W6HmI/5tsKa7PG8VDZ/798BdL96SPs2DsQ9UN0Tufe0LWu86sIKpGk4dgdoY25skizM/iN2u8Rbi
BescfhlRbh+pfMEIpC7BtMXi8Db1gUU4p0eIUqZ2FIlBe7UfPuEw6V4gsVD+IBDxP5mX2MoWOD+6
e0w0qUzd2v17eskG/B2KHFHLEpe9THJ2QGpcJ140Pq6YtGwsn4kJQZ5KGsDB0ghugTXTkw4U0HOM
KRVcarPDN4PIeMFUN+up2nHBCG0t8bmqJA6NsEsyKt1JIVi8U6Kl9jOHhUfs/F5+hEg2Jj8IwktQ
wrMmwsTizsmLjLQIa6aG9ALQ+YbkgFj45rRKmeemAGsEM1gkVg3daMDEWUryyR1FgfIjtTEtYLjq
93dGbl6EsZXcWsgkuvp6sIQBGcfCEz8h3+z8AVGN4uPfby+YoJctRqDWTkngF67lfx/9Jqkl8QSv
W02HswuZVvp7/r+kCsxYYLXPR9fu0PcxkgCyoM5GDvU79Ab6QoT6wzR7SyKwTSuXx5Fr5VQvIys8
G2hzLu2eiqOo5TGxverLEqXtvCS+BE95xlSby5c8M/+ld9YqIes/TKGe5ZeYK2pOqXmlscB7usuO
/nRONJxuU1UQBK6hiHCgLravhU93RRul7EYylO/5AonN5CavNETrLq2OK2r634pRxUGwJUNA31fS
TJCf1I8Cpi/3rxwIijWlbBO0isvtCiNk1pcoCsnQPr70yDqfoKI778OY4DXtO6ZgL5mZELiwcD1E
ry3OVI2bGHtiTYU5IrYOyV1WRNRfdqNXNbn/401NAIEOJpeYQSTfNbWqdjMf/y8mBBlilv5IJkOC
Un1XTOPVEJDXn9kYtfPt5lJOK/dxiHIAeJ1JhouIk4t0hESPPv/A/maBckdojQ/B+E92jjOZ0Psq
YOIJLb+Qv3wrPfQs1UDyUZne7fp7huRf7LANLRijpPOQF5hzmOyTzJKjduzkVuZujX+q8/oNpI4T
EwdhifLfS0f8emJM7YUx17ujUCNfL0opimJvujUL1sX7fwoWZNbx3mLgXZDvybQpBKuX7cp36hC5
+v6JJFQNq1vbFw+DZagbmg+3QN7eA9tc95mDZQTB3/rKYCa0ZNTgWZ6RKScOcyXOV2F8/gkcTZyV
IS/p3Gp2Bs9RNEpKvzTmT0PepKVgJ/zRgKYf+xwcLuLGrk/aH0XTXX9tDc6UCxKRUba2ofAgb/R6
w1U9215S4VXzioNFZwEV28Z5g/ukYUey99tBVl3huIRxhlLhZdohIxzfX9cnOf45KkrqIG3djTbp
7G+QrfiNxP6RbcGkmh31+vXbVlx8khpXS1vnLXSIyl2D7DMFi3NHkBn5sbwkBoDk6ohNzZi4YbiF
y9xtGCcZmmJiH3QDOJrCXMHXJh4ZJ/uMReHEiUTiWgyYHieAOdFXn9fJNgQ6OuVYg1NT/0r9CYAH
eVtlkbUXJCOCYmFFTN0yqSs0ZIvT5iRdYp4D8aN0aBovsqDimP3rYZk2TlD/OsoAVES1My85PGCv
g6fgS3xVYyLNaMCSLDpbqzMpfb9MobRePMSSTIoCaW9Dd4+q26e29Wh/z6tqRqv03z+bNrg0lkI0
N4wU7npos+Bb0ipCKIkc3O4mS9Yinx7fHP4tU2gGqQy0Cfdz33hTuVza30cbjzAWsVNWtVZPaLDM
HB+J0MGsh+T4Dyu0Gc5dhYz7o8peC60Rk6IpNjm/SUW+xNsvVYMVLTwpnG+J9H+GRG8E6vVZ+wwI
at/jvQf/hoD2x53S7Mv8QwNfBE51R9gSLvt+C6XffKlt7d02DguMxVlPH/dyYH5xTTQd8knIa2kC
CykrrQGUDsNG1fEtXh1yDoRRt8CsEwTmL2lfloVopZPThdiPZ8DlatZHT74T1ykkaFzQFpunI+Df
2a8l0C2kr3wc6K8lojX+XfRyQMDDBjP6FXT3eRNNcX69QNwrVP3YmUd+uR/7/xbMsqh5bA94L4iL
LjPNLx1d73lqVErZLiQ/xy2yJGPp2WB3K0Q1bf0N2hEklO15NratoeDP2oLwFYKBmByiNdF/VOaj
gPqv7Y7p36bcKLOQKgtP3kcBN8nbDjIt8YTpy1WfZ7EuURNNlsPCnDamD8/LiJD/EZI3CeU4rtvA
wpglXFZGiaFZBRFic3mxS0AzHBynwYALMXWkmkRfI7zZNUorX077+C5gpYt3vwNDCNdma6M3Twrv
UZCysG1yIvfQTBdbLFxWeA6SyHHOvM1Yy8uZ4PhEo48p8tMGOC4QR223AKuyBKemPRk7dARp96Bx
1zdd0Qt5BMM2zjD7LvQYvxhLXUX5KSMYjO0Bnc7uS7Vr6WmFMGHQyw8w4F4PNpnMfs3cDhaJo1Xt
6E8h5F/pzBk1zweSgJf8sHJXVF9N5r2mjmklvI+/mR+7DpM5lnPbKYfKdYdt89EiFktLd9LbXsX5
Tpn/FQjcdpVD86mpG66B8KGXXgqjXMGIYWs3IsLa7ekn/rUgpl4tmmXfFnFbOWUVDyka67EqEBgK
CIF//tdiFpLbK6NIvreKdIT0FF8kVSvDvAy/ZwCRyrdyTAaE/L86v12ngP+L88V83lQsEOUQmHdd
NM18sV9KlkTLo7ckUOk7INX8bOI/E1SdUleMTa6pBgOY0M35sjiXxxSmDEI+PyN3Me/nzwp/KmQa
yRANV7yLfYPiJ3WpIHs7Tr6NZr1aHB9yzzwp83xCk7yz95WjJcRejmZV/bMHLjZLJNjE/i65tFkI
7BbkOu6aD9Lh64fkTQM6qenYp25pPQxjG072deOEIIHGatCleTO8cAKhy72NZdpHGzKFHelHRGAC
hV+n9KvluzCIbiDKxZ45xhekqEeHrRsPzinsxR4aB7MycvD2TzlgOYdYmF2EriqX5dWNAtdyVW+f
CA1i6xD+7gcgq1YFNuIU5FP0xe5MSF2cm8JhfL/DoxVTuYqv+V/g5DBiLJwNg44gRLdWqbTMj1EA
hAEwNc8LhaHdVNl1gL/yIRTDaAdVYVHGLNMLqUoHGTi/qXE1CuyPNSGpYa9gMrRGql40sHW3iEIe
sEk8W2XZHXxNQgHVmd5CY8HzYfx6/np/VFIFNXw5w3DPGmysrX1PtLzh048iH9CQaU3viGBYIIOa
9PZxoQqA3UKx+UDirR4N+51f/rpqtWIhSKGPLuSdCk9SxzQkP1WyUEtxZ988YaEHznuuNXmd+N3M
jt14oSHq0xA8+3PNK7QFNb6albWeFbaHOGN4nBw4+T+BELWK/cd109W7lVofor9sdwIDU4ZXutCy
0g7EbI08wOBg9f5lKRUhYz799GZwpAqFuaIpevZm3hTJD5rzEoOJVNUYbOwZHlopyXjbG4dZiLHn
mU75bDDa+MRsw5jBfZnvdvTgkxdbRN37mJEdVLBCP4KlG1KbMVzAv1CJ//A2b/iu5dCIGvv/Z/MN
b4Z62uWLOp9jM8PU4oGlmLBRZio5CsHKtBx4qSj3klKsyE8sY49Rk5JDnOwfYShKKLmeXGSoVtJQ
Up9/moFi59XH+iiGbMl97azVEnT9q5A1TRMz7sezz/yaXSPXPYRNsZuHFsUX9DPYjNsx8D2Hy5A+
N2CnsnFXrq0wuxXEJqzp0McPRqypMxOdyIzy0TWdbKqfsvAzs4+HclCEykID6WBC6oRMKx5vwfdr
SX0a2g9fJNa3/28ukhPc5ycxfovu7AvrPYkjNKAOGGD5fpcYZd269982Eftla+0tHN28hAiTTPRf
/eL4sqBxTivhHXWStS5UgIoMfzfsMFBub2oyhLGVfMyQzuaIcHTe+v5nlXzCzndWrQlPO3gl9eg3
iFg=
`protect end_protected
