--
--Written by GowinSynthesis
--Product Version "GowinSynthesis V1.9.8.09 Education"
--Tue Apr 25 14:52:35 2023

--Source file index table:
--file0 "\/media/cod3r/2f2867b9-7e02-4998-978c-2568917571bd/Gowin/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\/media/cod3r/2f2867b9-7e02-4998-978c-2568917571bd/Gowin/ipcore/DVI_TX/data/rgb2dvi.vp"
`protect begin_protected
`protect version="2.1"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.1"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2021-10",key_method="rsa"
`protect key_block
Y12UjNacgHwFP8jRI1Y8NUUeUso0FBgzCzp9dHvMqeI/Lg/zhZcoc3McYPd93Ky3n+d6jqQDMwal
xhWVRJ67l+rAmbVDN2aNkoMQN7eAehBNBLtVQqvL31pMxfx5EPRIc41lwDg8DoCeKYeiegIZclJi
cJzbgPnOjIqTdLMdJCQjeQJ4ZTyQhk/1benE6vq7G3YtZdvKFnOMh404Q0rqZZMto6l+AVpx23e9
BAJmNSQABs4mgF+wpOhT6KuKXxDJCYgOG0o79QUDJFaKLCjnyAfF2l+ZlPFeV1n8CFgfsTQuvvYq
jo6B9HC9FoGGd0nRa4jYFrE373JYnh+gROUXcA==

`protect encoding=(enctype="base64", line_length=76, bytes=69408)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cbc"
`protect data_block
+6Xw8//X9WrYxGUqbRUuS8EnV36NXjYBq2FCyky+Cgl4pD39+Q22U287sM43GMJNxhM+emBReYkC
Zddfuc2otWmi1X9q9Vr0YV641t6JyJiw9gEYAM6H0mwa3qkkfCWq5YE/er4BT7bIKbmVFJth++Sk
2XbXPMuudh/6eHF7N/ADiXPuNxw+mnZOsh0yQ1wepfuhsamCsaT4DnTNtuytHntE9CEFTmkz/b/+
2meLp7lMgkx5Cc1XSd+GyG6kjucqFIwpNucoGumnGtD0SAma5LGj3CGwJcEG1KuePzmyI4kmQ7v1
PTP5VY3rqHYa427v5r/dv+6hQstoqjhticiGbhtJneiBdMsCE7AchSyubgGT4sQjNsVF+rmSkMfm
UU+B3V3tec49VS+e5Oj8rOG+vx23CtXEgLDZduXECQuKw7JfYGDpZ+7OlNWY9KDPW1CTIPZFkXLe
KsOQRUc24CuFz4mqajcRZFW5J1r8JrNq4LdIkuZGtFvg2QgvhCugq0Rx40c2x80AID7d7X0Mjg+o
HPEpIZMLV6o13zPz7Hmz6mM8hJDhauUnFlqt/5iXzrF8LTlTOIcYdXFXku1gHiqmx/eeLMacnN9n
OEZWIMSnnHrWJu5h2irL7xpE4FzCTpYi+2aJsJDeS+zHdXD3wZ/tCFD/juwzb5ssn2wzzGfDSUFh
QVb0vJhh1iHspvwGBa6YdtNKkeizOuKUhHDiRZQJHdgskVrJnq/ssQO0eoe04gBnMpVIc1QlykHs
wf6e3id83P1c79gR4hpqCakLh2VO7fgCcQs0H8E70Vb2cryLQ9SYwowo2mMJLf6Fr2Ve0HzqzhsC
fEd2n68kQ7GkL6dp/ES/0jG0NhRSTyIxzk4MCY+DHKKl/Kl0otZdcYIA7E07oETQY24uFOsSEdO0
3pqI/SN1Q/EYN9ddD6o/M2/IYYaFiCF4JbkosTK7pQdjOv7kHGNcI8TP3w0AvV6zq0wzcNPMK1/g
icLC2RVApSoDhB/GEMOLptpXiEi0To0yhNb9Y3gstGlWpP+WHejVe/Guh1UeVHkliivuoP5+WVvH
Msu0b6eYoOi6G+723kV5OK8VCb55mNgooxalBuhAfAFXFsNlbFqQiRuRkDmNzdB+joKFPhze6XQP
oCWgPOB31XPQymh9O0ldBpZbD4OhHjNoT4QL39xL+P6iR/RCdat7Kt13BElTV/dk1viH6CkWcvGI
NRQT6XmXfdqOXDK3V4VO5hWbRhE3WTayPyhH9Yrd256S8cdELsD0SvXj4HSJEhx6kf2OTTIgOpY2
T43MRpUDBbFRpXLP30Zk1OD8VnFW2HgS+JK+JZyJLRlrMvGvAW9+We7ZzyeMHqzcVBkAcYER9knB
eUfX9qlxr6uHKePdqRhZHADON3s8obEgxSguZzwvrnRoGhM4SXa0DKisRQ1rLVfGD56YWAcDNAzl
iy3W3X+IoPAdVmB3aT9TAUmNB2oesiqzPA/eX6XMLILYal+Z2bs4PrYVPj8p8t6IuiDKwMWoZyyG
jCYV+IvsXUmPCR1XPIeedLsgs4gK26DfKhm7m4Atn6OMntcKhGhgG/MsWvHR+QLfQgD73HQhGkaQ
c/cg9tHyGZoVwZ/nijf54cYdmdHCbrmv0LWZBfXuTOtJw2lPz1hBDUHfFhfw99HtXSi+NqA9peM1
Uhz9r/f8qUgR0K1p379R/sYGtxGv4JijDwAe3Fg+PNzo9Hh1xngceE86CqOB0gMvmJDrt6qsAcGE
gAbePDwaiyLlytXsFnMvbyPAILe+Ys/e62ZkKjJQO0KUxyK7SZ+0Kl4OGyXX2ftgwfuyFvwN6ORC
/6B+YsQxDkjuleqYXc9rqZDNhgZ0NU2S0YiDeTc5gnZWRUNhk2pyttCMWCvhjQNenSlSyNRD1y0Y
NG0A7ove6YdT0LPG2Sfqwg35n125vLM4cvPjJD7PbFoUbpj1cxCEZrASpDzTXCqa//4w7d5m8wmf
y1lOS3kAEJhGmxI8rOVFTfN721QSbFC4YCybkgTqDPmLM1SI3j6h594iBru0nTf65aQyLniqXk4p
qPvsgQGR04v9QWJGRWvI1bFsNPA/fJF/KXIHAdQzOuNRFXfKZsmEm9hWtMHOogVBbVStPuJmpIcY
hxGTOBjx8BUDMVMj/9Xyx54MrMlhu7+0V51qYObZOto4OO/69laYlVT6XdmfYcRAQH9wV/TDlx5l
l38kFRngMnLNYhQAxS+cSbI5ZFIb6FgzXv5k1Pft8/dS5tXubUz/ft+pIJ7+ljrNBugdq5z3alhM
N+PKirrMKLzMWIOdtzu9Hv87TOHiWmGZkQnvnJkVP6p9DAVQo2Xs0kB03sin92Sli9dNldr1u9Jq
+WMTQDlBGZZXeGu9XIjbZOR0xVAu4y3TNvYcYy5ykQmyVTcHOECGRD8JXmZ3Do9PX3ugKb3QwXZR
8H1+z3MbZ7Ww5MEwNihRIk0DtP0G9GaXgF4YTgsPEBPJe/y+r2YNku4j4IW4r06y9dKZ0rAT5KEC
0XIoihFL4jNka9gOBwAbW6nbAc0Z5Ty8OrPLAXG6K/xnDd0mgzkyNXPbueNXqVzJUy0U4mqevDfh
2cx7YZ0ZFhr2CvlP2/0ZchmCco8+HMF3Pa3PvbtyFznqc5eksEr0TP7adgriwjUZ2W0w5SOxEOvX
KtYKG+vLmN32Z/MTAnQ1yYsSKJCnK7zx41hSma0/TxuP6Ddtc+mC4IJGut3vrp+y+UE+vQl/rvzc
USdyOnIZy/Fw/J3KegubFyCu4UcgMDpCdz1pK0uC19gBjizJHZvA4VchRx3yaQGfq2TDg3wiwK9F
KE+1AuB3Q4k8XdZzgtXhtNoA7PE+T7QuE6TUVwmdQpCagCYs8LWrgvyCtWZy8tixRZbl9b616DWk
SmXP0htUZxlduRYePML3valU4iemb65+cccG/L3pwnI0vngcCAMe+NKGjPFngw95LKQrqxfdJ7+Y
XdE3X7bnZVOZyOY1eg14+1zfa8IurGBMhattnGYL7wDltoTy2jBwRcBed3iPtD7GgjPFA9mgO5LW
9IllWsN5eyr87+Mn167BsFAXtOf3U9Hjjg2t8mxIo9lsQemhjlsULNzJUjigZ2p9epHqdX8fFRwd
csQ+HLI7yo8LjVdTljezjBgHge+IlSpZ1GgJ3lPtBv5FbKkC/Y/U64mptnkRjmmdi9pZkZBczMOx
963Fm/qYA3HV090dSi94T18eNduPKjn8U1b2w8wogrBr4R8qPtyOEXysbYYkcgWBOHfFVTztYTqY
nU5BWxcnfBr9kxjO9eJ/RLd2yNIO50AIx1MbVyT8MjlhSEJShINwW9urBCWp9O/PLMnuMNLlKKYT
qhsmjYcCxwd2GQtOL6G+f5yuqwy4PUGBoXSqPF4zPijjDEZYoRnOsupESdpyDyjjfI7TLn3oIVVJ
5iglTIr7Nv4I5WJ/7LSBEw8/bjyf+0mOcP/JHueKIW9FVW3Kt+XfwhvTZazI6YqQIAZz1F0fHKEC
01rcvAJslyguaGu2G9UPAb67Ha2dUhAOENB56PxjYeqiaVegtYRpT9JzmE2bxLji3NVHvIBDfUMb
AVe+rJyGaqdoSo0ZPw2IR8gGiot5BjcZhb1PAm7yta70V7AeD7095SU3eCsW/oXzf3q0c/b07FGI
+N5v+npGkvSyLz3nKGoeSknqDKknk4EYsYL97BYKupLwjOzg6xxBzpUTliwHAtAg70oUuxJPOJ2J
YvHhxNcCxxcKH0v4Gh9J/+FTo/fmG0IpinZV5C5j6QYaYPKTse0YZs/IAO823cDceD8UNmmjYoXK
stlBqX9z1xaWA5VoujQ0k40pDRqizVBIFih5wiCbrplaSD9Ha8byQshFsPh0LTn5NApPmA0M3eRA
dhZ2b9HVWT4g8ddS+4TjZHoEOEOFtYQycXEcJe0uF9sRo4ccY690wNfZ6qUzJPGoyWNxVzznGZMn
VpAEf+pe03s/3pbS+3lFweom8EjFeEFi2SP1Sb+uHswSrg8FXYX4PCYh7vsg+rXp8M6EeixyPFJr
bC/pQ85K8ZkxPJCxm9ueZoyOoxC9zQi92hd5kDSJGMZv9WnvL+EYwZQ+3gSpAju8OWeU1o8Y9lTw
WYLB979oSJNo5jVmrKP2RcCWF+Bvs+qd5CKCazH8Hym2WyPBQiUZzwypXtuTccHRBA7EFC8l5zCf
Jc8BPBGxzFAjYmKfCiaX/okL752o9JQ9iUXkhiixfQkOglunZZVMnzUeuMh60RjdevE1Yt7wNcx4
IeX7LMc/2d3tS/qU+4EoZINvEfbckK57nmhj97AdGC1tAhrEn22lDzmBvzRbC7NeGKPP5oD5hXRM
i8dnMHuWPC16UyKkQNYh8JD+00pXquVoMGys/WgDmW2GY4rQm2qBWyl7Cg98egkEj9XWI9TMugRY
Xd9D5guK+VkbpqEjHee9ltQGsCoPZlyug76lybfyIfBwZxFNJokBhaNeix4M+JoaV5WeIIqJtqrT
Y8a+bysrk9k1gAnv/eF6KlPrxPbGs0Ft/JaABQ4cioOgayFu/Qtx/ibWh9GKewDShNIzBrZLKxiD
Ns7IWYpD0WpzXRuFmxZjFYoKFd+bcbg7fhk8El7lfvZZJMEDpCpAwgrpQQKPeGn2dqVjkQ1W6dVU
+6Onts5mNQ9J6NXRXvsGyVJstnulaKfu2+1g14irM1I/zxlXPvF5AyVJ2TotentSKUC1REvGz8iB
QSB84wie3BcqPLpBvugpAwNruUQHCEZgBvfLmOqgmnjY8UYeVSyWl3VkntB0m/PHbn78VkA2GyMr
WtJzF7RjwTqiMKm0kv897EVZxdNoQ9HxgsAeDgY7vfFrkcx53q8ViO2DYS/VZ4aQy4/eSDSFffvg
dKkOFXKk9j2k42NBFubFSYO1Y4KXaNbgwnp/4R7Drfkh1Ui1TfNxDOxY8s5h4VCI3fiIWHpCOJcQ
dr+Ts/9JLE00MNq84Dq+Aqz0xmvRbXZuccMwy0Qsnt8xdcGJgnGcV4R7S8jopqqDpq7tzBUqd33C
wSSMmoAsL+bBpR6sMwDPzpXm4K1Or/wfPZSjU3lUvhCVXbfqZxsUkWWYLpgTje+e5ExpOWy10r8k
yJEJBhsa+MMOwJDVM7tMpwoWwqQazNHWBfJ5biAZ7WVQqZCAbNlKvQL4TIPKY2JXxj+3bMWDU9V6
195BMSlwAHdMk92xMJlqtZzexYEvpItZUVqklJ6GxXdKzFx7r5T/otjvJYmXCIjabXQnLTYZjQo2
+hOb7nUNUMdwComUZrmRcV0L/4eegnOop9gbQ3pjBEGRRCL6fhIhefOBx13/xmq3KQp4YKVgsK6K
eV8w5SH7A1ka4RM+GLT7QLg0kfZU1GrxhxU8ZHyb3p3ounGHOaMHy0O0tS31PgZy11bqhdSTFKCM
JyaDH+lmuF6W4g58TFFMeC67r+LAmq6WVxT1ZOEe0xdJS5VPLTHJ2hwNWvFnrzNmbtKwAfl+O50t
ZRT5sPP0aGP25cs8cMBhHq07pGav7bEgu3DQ4TuzbI0xaZIfyPYdSs2P/iHpdfqrU8lv+3nE1IKs
3BffpP7A6AiGagEAXh/SOQaKkJz8ekXNZkz6Gux35fn7RdJmfMCEhMzFNca5FvGvTy0QEznhNLRO
4h8uUWWmioY/XVhZSMzgCLvCGxZJ2URJkREAys1KNEfZcbPfFnE6zYxImCotHe+ciUUvkWm2gAl/
KWFlLP471MjDek/duDsnUm1qPpxxJVhvRZ5o0h3L7UhYX4PtCsxEHZMPPAe5WJWYOrDgHNLpkfQb
T7Mf0sR9zO3lCxrOUJ0DqZX/lD0AoASZMg/jYwYFaN996sbCYjpvqXkleKQfhlDwaUIPvgB7bTeK
JshUALM8aZwtIPc4wkz4rHDEBqq2ZCkqbksdy82MX8YSQdmyFx28Isv6r2MfJh2oA00cNlaXA+0B
GS11320FLcgLooN36HkHjmWQnjRSrvZs0GnMOB4UhRKzwrWc95BWL4O/omcs6yTK2T458YRAmru4
9dJJM/gzLT3phQBUJv8/EjS8kPBRZB2kfmIW5q4uS6ptaLgONtj82ZIGb6n8p9GMlQi2Z9Df3R3j
g0HHaoAs/924+FisIFBtxl7zPTPHOTFA5ZGoxHdSFgOCjPbcvcFZOmhEuYYkyN4/krCrZCO93rt6
O8JzGgvRy6+qrX/n6dLUPAU5ckJ4SFAo7Y2SsuCXRsC15hkiTmTXP9mNVg5vtVw2Qy15pEjKvsTR
vfM8EQPsb5BbVC/PZkUx26CuMN+GB7FtKAS913jXV+qdYubZR4n4WRfbn7tLBuZItWbv2rlwFA9o
Q0MBtY/2dSu15S5Mr6jWfr2QgZadCv0gHQLadXFTft6k3pZC/NrByFfUjiWR2fPzZXOM69B/F9nx
DxbPhksbE8foli3CAxEKLbyMt9FHLmgy6TbiLWf55Co4S6WaN+QT6haNb3fLpI5wb+6sYboXkHbW
K33u/h3hT8uO6NbWgcIovsQUN7YUD/OfbeYNLReA5ZFfVhFfx9uCYMyp+8w8JaFf+cyvE22aGvK2
AyY3/pnJmYVHBEFRqnSs6ZpYY9S87rjyKo2KB0gVWxPa9qU/VpNjurTti+exf1n8nwl9i7CzSBLA
gsgUW4vBvuYLldl/esWsReEO0O8N0VfM1hbfDMFjyskN6pYb/Vr6cBmcip2b5BmQ8kUWDAJuABKX
byt0LpE+UQNYZeSdh3ufiQ8VmMskBqV+lS04PObihSygtJyvqT+PMhdI3ZgKzcIjmy8Pu1zagfDi
OJU4b6sElqYC+WLXjaYQcixYxXa/JTr8o3M6BpHJ/4J0p4PhQrdznv7kPE3aBnyQW86KLaQVz2sS
UUHzkMP9PQ4InhDofiu10U7eVf+Gn+G7G3zwCJai0D/XaXupbjVliB3d4yZ0SzNzrBUmx8c0zbYl
o0veRGrh1Y2vi9P4iwXFXqXyLVue5/K8JlPbRWSNnoKfqurzbv3w4m+f/unENr7EOUUOHQgCOoE2
tJnMbwF70yes/bAp2HHWnDPe3l2xfovbJkb1KY0GMIia50Y+jeIYRNMZSpmaGRD/1dRP4SOM56Up
Re2VkcLybmUQhAnzuVMk4epLZ4Cer2RAGRLQ5Jm0C4S80KtnyRLpvfq86/VYyvxzs/WPTf1cVFDf
J0ujVsp6Vfmf2uQ2Gemr1pu5iXJ8ZKylJtLOu/nHNnpHgCuJ03qHAKH72beykhWSe82L7zXVph/H
KQYY/6UgVX2QqqmCY9sRhmrTJXKWhF+z0Rk133zBhUTfWK3H3ibdjppOtIz0N+psi24Q99xKmbll
EvyT3mjzEarqy8B3zRjBkQ+KKL5Ya7zbJExZfvX0GSDGsy7APP69ZoWRC2FnsP29vC2iDNITtQaI
KcersdzhPzCt5UTvwA90oPv5tAtXJiOp/4nxbJkODU5ZDs9OyO4DjdMRYwNWpI/pDAfCmK5ZteT1
L8pHh5FE8FCWnxgrthXTpB/FOC8DWjEqfjC6aQvAkk68c2Nz2aa69+mvlJa/beHDYmTUlIhx3NTA
LnQ1wMS1KezX4b35EtNBC4ONngmCSU69ovcjRsqj/YW631hEg3nwptIHOvbByulM5Jjn6Dhqmz27
9Qj7sS92UwRUCsd2PvkF+as9iMBqxW/i6h0Z3sVd+4YCygeRYGdUF1fMwJEx1zPRqB5piQUshp+j
TZ84dWO4kgmU1UGPTZxe+bNf0dlYWQUhq9erGhZD6iHbBSGq6eHcdWphl1OTDVQmUxV63yrHO1ue
xnlxw7zV+OUjtDxVZ5+3dlxHZ+9lscfZCUHnMa8HGj+crS42LOftfSPY8GC30G4JM7pJtzFtmweN
2/dG/QniY+McwqlnewREex4HwXDLWevYhUuSlDAKb0O/+uxIFF0VDCKwxXFNuNYRcEH/wVtaukjk
8+FnH6aJp5CxcQdSZbcdSSR1Ezcj4Ru4FQ24T9O8lxGvy6lbkixirFKfYYCMT27rkl6KKZKTaqtE
EsXSYvtNagNsOArIfzbM9PuTyNwZG11R5HV3mUq2lHpQvwNpaHZZlujZ0STJRGw5fWK6+ZDtqkf4
tBScTJ2scuIRj0ftyuxf0/sKrxqjd/zdzm63UN1vFH3H23IERLOFyV+6vUZecsuXxzqsSys+tLDK
RVfUEJ5wXcaPKI/hlfnWZUTuGgmVxUEOnlaCt4he9bCB3sXHG0T/0KDhxFIGXLNKMOQmiP7iNkC+
9noJwV/WrVKYkcayGwicR+cz+LX09B0TvSpGTVBpnTjlafX2Ahjmm25Yevnig3E5j97Xu+ETZV4P
lmrR2368KxWGX5whSKgJncxQuK5PJN5cCulICNimc9Db56ORNjMEJ6HQrM+vpCWzVHHD/jRjlJVx
+xAltentQUarMgjzpawc08Dy79qJMYFxT2fday8zXg8ZYS0TCX/wKr4EWQu567aF78YQB1A9jl/F
MSoRUfeBy8Gg/LFaEe4AinvBdOJ1ov3gHi63TCcP1US6UbCQlzt7ubzxLO1WbttH+VuwLe+GVnJR
KEIK7T5ofAlwNp5lfJmfBRxV+qEQHkitvlAfdpO8V4JyzF26SLz0YBo6HeuHmRc55ZaysJpdsIPL
XCq9IRKOWW+nfeYY786dyqTgL1YBor5iCeykT9YiSolcLGBv9vTgUa+qZM/wPHXk11XFbHpoPJmY
Wck+8C+U+ERNVfJqcMnsquzB9cDehXE/DyBNL6foZvkqvaAL2rFS+BkjWrm0WpYsKerHyJMlqbr7
r7diMfk/sSDsTiaMbdCfUqM0yjJGv24+SkyBlIQE5VKk3N/xxAl9RDtqbc1pSkxGHhzHXDtH1s74
b9kt7X+lnCYEA33Rjh+EdT6PF5DDR8xPQLbpPKUDzFBfahqU1M4U/d8r2nLWazfQqVM24mAKNO7r
18k4z/ddeV3/zw92hPBfLmCla3CirKAIPuNMlFve+YmQYjY6R3l/T5qIyNVwgiIJIN34GwDG87Gk
tVg/ZR5sKX8EmewB6SURKky2SEkro7vGwHCXGYb/l2wc7z5mSw47KnGnHklXXJTdgsP27fC2AH6O
kIh8JeVTscab1nKCmV2tZaHgTn/SdG8COh74q7YsiGgbVVauFTV0P/6HYu5EjHBITcb9XydCBHVX
83zZxYEEx+QJSVPBpmGYunm2Y0qrLLUsOt8mrYN/XQqXfHdwJ16DPNYQRrK9H2LeNpg2d0sQo1Yi
WteB036Rlo+lOgfOBi/6FisYvhQTLpQMKHVFdBSH+xfR9TvbEYEP3nPPMqcZHfMlfoJMpYUpfy6t
ic0I0gzMOG1U1Gdv5bMRICNGk5/MS9/j4qkf/LR7fbOD6P2tC/YyRrckiE1DPRBf+CBSepP7ZuCe
VCwJtyzDI8HAQbZZyO5tWUDkCup24qrk65jR3alCZX0T2/v3xAw047T+GyPnpRP/STAhNQgcyLdZ
O9ZzEGy/PwoaEw2F4s5vLMqMEPeU0RV/T0IUYmd24fx+Kh/i9rVm9/belWeWLC1kIGa7qu+Cjn7o
MVzgwZ+ZixWl9oPw+zz1sGligzMOXmwor51Vsn2p+Lv/rxUc+uYmI/aZfK8lTkwx4WlEOPAJOvJM
DDD8fOi4YwDSQ11Ujr/vEy6LNNmvzWHX+LsT3eiBAaz7+caft69NCrmfyNQ749Jo4HTJCO7Wztxx
5iqGVZdT8q0NyXfNYAFmeq557Ixy97Wkm6U6LT39c4cAsj2h3VLZ3zW0Fyn7Y8xXok0knZWK8xYP
9P72CZTbYZ9Iq41szHxjiQ09TZZ8PNwt6BD50vxYznY3be7L3OeZoXs2UFCLKn2nviE+ktZXmoR0
PJmI50OrI0tXT5lVIbeZR7Pt/1EUar9vXNzS5n7TwFZiLLSr6MUqMSEQA/N1rcI1dVLHuwtEqdg8
++sZFfbroCWfeGeh+GoGpYctbGkmMSRzvVRn6MBtJqSrsjC7e7jQbrPDV2m21DQDPCcYxWCTMxI9
aHzjLJLPN0CZT3fo8M6m1raS1TFgsmPGXdwqjZ8oSC2iaoCuLqPvTaFAz0AHXb98JmolQo31LzLm
aC2Ei3DVOmC4ZUnR8nptnzITWg9ryPouZSDvU7mKXw2rpYre1HKHJv7R3OFqNPP+3QCH0vcGPZBQ
ETZUecjmCIj1EKVAtq/AjenM3uXM0CIi/GfVdrAog4YjHYh41ThKGiCD+F5I4YD3ILEhg1UWExUo
U00ztsQwRUyLEv06c8R3kLNcWC/uBE+TwDu4VNOu37MkAX4mv7JKlDPSwgp8bUYot3QthXV3+Ncn
v4zpvmvH+ezGonJIV48XreCyUI15BO/ZpYXX5TP5BgW+ESy7k76j4DZbIWPaDJgsNNIKZGcP6MDj
6LSZexisqPZeCQVs8Wo6VxYFBybT6gYxhl17cUTyFFSnLLAhzsR8sdJwEk1xu5hw6acVp+fXyKXa
Ycz0c42hdHwPUg9kIXGzkWL8wM8AXjeG1ctK2o4ps3564RLQhs/+NoOrCOkOS0obtP6RtSLDyVPW
ERHZ3XlDWgGIKgC1sB9Nv53em5pwJg0iK8JHCjELzIzr2MRlVEumm8Dhzhw1KDqmXz3cMJ8j4kgY
hBRfmcuyQ2V1jYS8+KI11pWm6XJO/WGJEWct6ZnHAnmtxm3dJ+x6lwsNF+UTfFMQPG3C1SNjkNK0
VAz3C8Jgkq0VUMd8PhIifUIitQXKBpn7WTZyrnNXTp9g1WTu+FwF2Ms4znBHoFuQ0EMPZFxz3gE/
HqZEFuiTY9Zo6ZBsBJE/pKBcruVu8hoFHF2qa8IpIGt4lyOESMBrXJn3pK82pMjM9qsVPsTabkua
pXIE+rIKyvcyZGaCZ8w6DsdUMNXXNPJY69oKhMqCIKSPGQvwZ1OcwMAfGrFxp5Qflfcx7SocCcz+
co6tgqhlzcmzBpR3RvwEuX7ysemLEERSEkA6krAVxuBvCVMJ+eRq65Ejm4GbfmIg//fcZFB1zOxm
YcVM1Ab2jtnQZsg/XjnR7g6AEier339FXHJOLU6fyDaG2eFNP1J68o+Qz9IBl/V/Vnh/2dkMqKk7
chy0j4zrEE1SMBSo1HByS98M+gozMM/59ELhofYhoYr9vxvOwDMjN1czhxPdBNYgqUTDOx6LzcIG
fAxLJMVhDYK8UADGzTLMrFrIKV8mPpr0O/BFKoUeLDA5m47jpSIqLcloQTx7mbiRDdJg1Af+LL6t
BGGXSkUkjpkER5NieO4aNIj2eAAJg+rTjfGdrHdILxzrPZnV8uL4scpMiXSazhQprscXxL53T3Tv
HvvWGNTtjZ3F93ttIT203+YDDRhobylWhnsmSUGHqXsJRy8LEHnDzngW3FTrMMmpUT1oCug5PuLO
vTXdBF4Hg0QZyZD9rq4+AOQwpMX3dQNzxDvx+eJaNjiZnTypz09VLqrpImYEa736pXBBAsDxVPkz
kDEDy0BbSBQjPTNAXkWvHc+T/cskw/UMaoggVP2qfzXWLiuPBvqGeuJgEvA51bwlQa2X9yIFunTc
zS62eZkTAY5zulrA4IRGxUPONO8x4Tjbxl9PdWa028mDiySZubowdkDLGEHSjY5izvWplbKFHFDA
ewrzFgTZ1YpOsIzIwIWzlX//zzW509t8WK/mBBqeN+Xfgh6nmRHK6LuHPVELF5el8giHLIRJ8bUL
GDAcJwDkJCjV4WrWTEaqJvCjKGAzxvtFYr4ib9ZLrcJUQ2Cmu+0BV1hfVYB5xTmfYlfrxhWbW3JX
jM/k/5XIrRHkuQ68ZHtuVEFswOoAFDnVaGBP6/1HSom8gL2sWrUT7hTzsCwcvHHHjzuTgzM5sqre
GGSPSV5eOaQslE0Vfe2B610oXD8dSzqg14DDKtZQPhLN5RAI9SRJ9SK2KE0JqYoKS9gCeovr1khw
lWBYLRX60GJH1LSsEI3RyWeICg9aNYh97LHxQKUX0xJOJErkSiyn0hRzMYRHIBXqiLEE6xFszGMU
7Kqqv2C5suBXSZzZPbl0B3xIj3s9Dr8LBGFwvjWr/5II6dUMJrls0DSNCvbYC1BZoRCJYfZxSIPg
WuqllgeHW5oNTz2dokiSOC3Ynl66gU8scZp5Ds6TdBjf6/2X86MjVLLxkiRxY3Y1kW+cCg4P6N9U
nSZUp6GTjTFqze9Q8BEO1OlIwVen7Z67Bi0zlDipxkGckQ8j+CYOpmCgOQmaqSjAhugtX3d4268e
yrWMN/2oLzyi7rqyoklPXojWs74uFeA68XPjj0mDRox6VkjBGzinPuepODtCT9DbX6sd3cLc3DaE
TBiznprYIYaEhzdsxL5sP9BaLNvd25NElQfM5LBULb4QiaABu9NkTl9nacfcQUwpNuAkpWiID7E9
Vbenj5bToPFCrkF6yOCOO6u8GGxCawim/NrIGWTZ8E0pV5s6LEkFWsWTM7Vvs+FX/ry7O0mD7zxE
8cmIu7BeFivhXcHLSmzooZIH7QjASZYFunwAmVKcAALjBK99aaT3DMIZu+eC7IkXoEAUlYYZs9TF
UCNMXOzW8fmMzmWc06QVydGg08ZZGe05p1yMkzSi/D48U0lC1xQe3e8VecMQxrKGi9wqEPohMGcl
bpO1VlU7Ahd0nOralc3yviJxoOq8VmG6lFYDdjusW2UxNgK8smmMiLq0jsNFLi5pFYE8OICnlLbe
RC7s4NDTpRqbUXkdqXH0YsytkgEVKs9imeOU2yro0G3NnbNZKwa9JdBXnMJp6QJJABFPevLX0hSn
ESVKRj/hIIZuWlnoTtuuHwmOyN+BkG/qKpwPgR3YDIlyx9bBbzODeg01DNAh8fpH3arDzkRoEesQ
HD8ZOL8N3o/PLBgNRVltaicLS+imyyLFk2QJRCQWqSHnqYM70+BqCJz136pgNC2fxZHY42bcGMDq
OnS6hc+GMKGDgWoPtmD4J7GvVClrc1ditjfsOmzRI48qBWP9CTzePpS6ob8o36vFZGU57qtuDrQS
9sPDFS5rxeOtGt6VaK74u/T84hHxFewmRkSo2K98Mz7N/0KxkXXzlOF0K8nRohFBBME3kYfZDIFx
GnbM6ayRpIW+VyQj5Lv9PmgxYGaLsuyaCnDCo6uPBJfeZv0BXQ7mfXXA7fTmbTIO8xpOgTKJUDZi
6vLuavguZJeRZasuyzNvXEiPnbSpZhEV2mJDLgCipV3MJBMrQqgOHDNK5/xcPlBDD/zBEI2uG/rC
0YAEIwAdWiM8JdW9ZDTP0Vl3rLpYBoBbq4fe+l3ClaMHzjg8xqs6mE5ebjUY9tU80sV1nAg+Ujsw
QHOlMrvEr7MyUADdHzCHwBGdtm48c93oc0dh1Gyj/3iYihL0WbKG84ky20w4SJnJaALEwgNl5kDs
E+b0/zXWi9WL9XjaVamY4CBp0GPkLGD3nT6gZ2Y3rauesoAoiaYkL8VyNvJAKCd5NqRdooK8vX6g
Xg9h3CYX84UecFY282pvACwwpMv2JYohqerVbnV0nxVZg5oSK5cjLg1yvF7Q5ycXYUaw0fS4+DP0
V1Vj0HQS1+5jINlkiV2Sd8XERgT3MdMivlt9ufLb18/1PLcd9FnJbaQCvIgszxFcoVtyT/ErDks2
Lf4DPRBty7NTliBIsU4U1bSioWbex8zO/5hMXwXZir49MCyY73wM8sssKEaFO6DnBdDbqWSENWEV
+9ZI8tt2qlLTGltftKp2XmxWnY/b3+cAjbzUpwA8O3LHpJibcX85w1A+AhnIiBmq41b/GezlLXmG
ns9Ror5KvDsXg8X5MxDeclmnuASbZ/1aX2iVkzV8UdOYfxS06U5xO4ABDVJRu6kSRIzejflF5iiU
tEKc2YkgKbUvuznmA8lIAgQsRCLx1HiB2Bv8LMkZSUgWrnHNnUwcmN2+KC1Hz7/a21qoaCRxyOag
DU7lIRti0HTSM8GPWfUEnn4DHu2KzzU/3PO66tA8zBAeV6j897EidvzTq387eMHJ3pudyoRACmrB
7ebzf6IkYtm9TUlKvgd3wyM7Lw5kR0E84yPcEccYNkcfjHkMNhSgqH7uCYo6+YdhiB9l6OeBFORL
9tudMqcIO1UVAK6SRExmAECFo8SOkh26c1vwwkx/zHIo8+ZYMmIKoV+fyzEo6a15PvHcP2rF7UTu
7TPau0pgL3Cu/SqWzB/jO6SSi8kP+JeELbMna8S84d0sBxxR/DPeqfhp2gpliRmjSwKfa117VPc3
IDh+dJUt+YfgUUfpqCKXqOCToO/MHaWjUaOAqaGxsHQOeCMWDKOSlxiO2HAyhhrJ3EEbMD0rwqZA
LQhqABAmRs92c0WL+D4RQNjbNpd/Qx/GrVRw5r7NjezaEZamT74sRcBNpszwJnJKqpDwsbXk4EXd
hwhjPANuCWm4Y37T0e2Qv+xmoKXtZ7qii2U8JQx4Z9SWM9XP5+Ted5tFtOatREork/dbm8+KeRDV
TlZrDibn15DG7va1YpxAEYtLa5EG7+cPRHFtQgdAp1eqZrTqFStbBctbR2H2sdeifMDWq4qFJFIs
+ALPhMxcH9LVYdbG+65AlgpLlovo9EZpJOD7+2aDIA2D5WCesZNVDx9roT33/HwOHP+01kCuSHMC
aR0UmJip0RFTnUinaCipwH2AiEgMgJz6gszVLYID1hwHXWkJtwvlRXRtzjzv7WBuh5Fz8OQV/gHd
pEyYy4V3dQwzpX4WRSpVQkN+iSYxbaIABIZke101HYlcSra7OnRZnUMqmDgSvFPlvGTdH+w+KfjQ
eieyObcDxYgE4NPD2kp3PIEZJQjtu3vAVXoqaMe6KvKaOuvwvOdiEvtU4VZsjNwnK7S4cAXJfMJG
gjk54ldeLHBNFyUd7UBex43P6CshnMQZhrYLns7IecC5dmEdymYPS9qyEgx9B6JjoXxNpX7aa8V2
hc1SV57rGQkuVjQ2IEuJDPHggsyJm7c/iaMSC9Zw0N7LtJuTYO/ZhMZAF1BNIR6WZZbI5T333l2R
D2BJkzd7c1Pl5lJg1cF0ZioiYS0SfaYN5kE5sbApb7/HBbTFlcq3qXgFoN48ay7zGS3IsgpbHo3/
B8FGG7EUqIIylW0HYStIFdJaEk7eun9DR+wqW5V3sa7o4fxPr5tfIPPnJmksTSH2jcDDDJtit0Y+
DYhX2ir4CbGGQ7M5riEEJsXINvVJHE7B3OOEmkxse/dlEoKWsTRMqVvyWZJi0wvSIzQVAn4w0pJP
Xff0Vg6NtW+UERgnxNX6DUB7RP3dYlJNO+prNvgVTrc+yuGZfPRnTPVcPuyWdzEUynG7mhb65hcs
mzvAzLW35FgDmkjqZjoqskXYp+cv6dnzOplhxSHm6itTlQTXfbKX523sM7DaYGuN7OOU8qbT6o6D
gjbNy7gtRGekLhGi7WENyxiq688RtBkrFjRe6SUL8LRWXkcrNrcu3RhU5qiswUDZFCh6/+Cs+Oqj
ay1/skwI68oeqdDIrp3X+qqLuW3K1ZKAtfYSTOiZ6tlDsk8OWBNTjbF6G0wrlA9utoqhE8IlqEEJ
WM25jnrZpNnRcf2pDUdUZ8tGACabzPMxmCoO/s+QAUSCi7oft/aFHvYrwr2Lf0wkqb4bB5dhVKYH
Gjx3C+0uC3UNqcm5ow1nN88Vv+pajYNFvYgBqEuRHhDz8CKbZwngURaRqf+SQZrqksUqOTbYNESU
DYiOwJSsRdxc+jzah/HGxABr8D9xoSTR0vL4efHRTJ0fs+KfXsRGG9Wx2FvyjDVLXVJkR0puoSFj
C2ofY9hxJIS81yfiRbuvqj/n+0glmO478maQk58H1ehHuDN/gViP18tzDxz4/y893QwOiHJap8+M
/vaJDBBQoT5ynkYpOCE6eqK0w828rahhV3KJ6CELCUUDKwV0Ey8Kd0d8ED6ZwzuImk4uq303KooF
ChrkMV13LE2ziK5os6KAdothvujLpWMiBMhLSNln3AHAtpt+yyfYOfo200HuY3yBm5Xh0Xd/v651
jO3HVodTTDcTkKQWy305iieGZ721yJRkJVmbA2LgEO498jZ28+s0+Xyv4cKCK+pqu0uS0e86dM7z
bVATZT8LPrCSQI29kG2y2HI8Of0MmkUqZkR66HF69RKhNEEQ5uTM1a2qURz+u1WIPdgrwh+1sFyS
Rt7Sq3Yot6TRoctcdTkhdMEghv8SAhJoJetk/+M+ffSmHAFsz9IGEWWswhUx1kaHq1ykIopCysjY
1ErSIE2izPW069B+XnTPA8jftdXtiZCvI4lPYK4eStIyiD5BCeoes1Y2OpSTgp/A+WXyoMGdggMZ
4qe0QAnfJ1fsdm29zVzMJLNrwDtVKKWMWAlIcbNqfZ0oCSviR+ZSecs9scGwIHAapboejxERwUej
lTM1ya3vZS1/jZg6LTb9h1rw8S+IkRSoxuf+y5kjLxKY2rmU0SXLk0H9pJLzVKWiLaRKV2518oWF
zoQhU5YJYAjIECMgQZNwPvjXinDDTU7WNoa7B+aDCnVjG6r6VyiaKt2JpDsWMSBG5yfAggond2Z+
bVX0u51fHyRAxllJJ/qrTLFBR2JVivumCGvtmsMDy6RgUUP+sCsY0GsiwaS19AMbTR5CsvlcOngF
fXy94qwHpCKKwvx/FH/LrsYX53YqNQygoWm6yK0CWO0y7vTNEAjBsa91hdtVrLGPP245a6YKFmFV
yBvxCE8PV9AHUPxg9qYQicg8BFposqoWtY49jX32HeUC5RptLF9lbVZ4PgK78ncL2Y7KnUJFRZoC
vjsIIlV94aQGImpjKxHMme7IfFPvzv/JHspDxtv01CVuLL/wfSlrmUMKzS5T44Qq2SPEh5jGqEet
xf9ZyVf27kW2MvQSEk1i6YdsolxrgE1S0YW6F1BY/49/AfFP7bg5GEJHK7o7LoJYysfPnhQZoOQv
+nQlOEEH9Ar0XZi3fRa73L2O9OCaMxjwo1LCJzhVmiZYyLfbqDw+CJuXIc78lnd+DcgZbuwdhY3T
/KiHnjtmIOMZMmvHvrieIvqkjeuraM5piWv9syaIwm+rm3FhbTLUjYKB/1E5bXBnYtbJiTvOohhj
+0ZoiJw21Ei38vpAvOebryYZym3gubLfeAd4983t7M8p0INUt8ld7AT4Eg79DqTJW+5ClDck9dOy
5MJ9Vx6zsRgDQRtsdFaYcUsWY8iKYiJ8gZt9Zey2h0b0RaZid7P5sKOuco5sBrtgCq/bWW7rIElk
8xXeCfk2ngPNtsyp++eyHjIVDmFvxXy1gKqqO903SafPb8wOVeV1bEKjg7U69eBYc5roeDXZuLh7
fbvjTsx3L+MDw5cSAcwabuWJwqQ4amVpWxXtzjWq4IHFDrakbUTTKJfMlJsPouHjYcYUL2qur4QI
ngXCbtvLcD3iRwpq3hsYB124GihD/BhT3NupTV3Pv0ilGdZMRnn1acmMOMOP7cv/I7qzPBhypv/r
5EV2lMfpvzSUykVmzS3iR/CQVd7y2ptxxrRD7lNjzn4iV0+oix/MSFENkHcaj1yywmPhaIjBHW3m
h7a+gc3JTJOlolJdYA+zjdtri3JsBES3iZxBtzRecTU5MFeJNmoTEmskYhx+qmV2TC1GChrdueij
gMNzVc2hzJYCrY9YOZyazfkZLW6yUqkBroEnMn/MKU/AqQtyHOvgbAvZ/P0lZ3b/cSfkfaIYZx2S
2pU8wHc/Ps2puqjVJhu/sGAyWFM5cfoeuCRXW3Rh6lYtf2Ka7VX+rhe+xkEut68ju0gVBISN/TDX
jRzeU/+gIc6Bd5tuyqUYDKsoP515J5sl/JX/GRGbzwsajKmVqAUbg17BQs9R8yyDc32q5Q2B9/l0
ofcWIJdIDCz9ZYJpYsCG/Ot3qwPukPZVmduIobWUXMjIxec0z4se2DJVIoS0cirlAkcqT0nmzFrq
UecTJ+39SxK/OhzFjcRbngtF875oV0HGBXNU2mrVXwjk2hs3ZRpz6LHksDohnwWQFfBKoRoZmp82
XVPX445FRH2yJgAe/8DAye9ZJUi6CvMT0t+jumM2ctBwn9gDIR3LBwGl+ztIEVZuI3xKpzszAX7j
tinFZLZ06c+skMyk4UABvUPvZd2zROqznzfDQInqggufMXN7Bcuh79iNmej0oV1yNajmMKU9OzqO
SnSXFvIs54oMhYrXE1YAsGH1mxTAL6dYKzXiTeSG7gO3oxp+M/+xzVESHZAbtzLvK9AzkU7++uQb
qzZjiPwhDxgNg7kRnCZ9JKDlLqoF9z8R7Z4DQm1YES1jqxSuZOsQ8ObnplfnhYVa8IJV3UsHveKw
3qfCkIdjq9/mBkvgS0P5Ku6GLzdKOI3F9h89+dZmi5Zz5d+xy9Q2jg/RaEH4b/sPXVNNylrZ+kkN
4Na76eUe0RsdS2Ak9dbQwoGE9pTHI351vS5JRgISWVwCj5hYN3xMQtQSmFBSNa2RanhCEZOdNCH/
Kh/QkUNORBaADZy71ZC/5nIGytOOs/LX4qXpnw+MuVP3OAMMQptwaGMgdM+IUfAUgJTjFihtONh+
GHC1UmPu2e95diimRvYu8xXfMsVnULR1LAbUz7bbW92Rz+5qewaSMxLYqNCus06gP423k12TYxuz
Wt7yuCPo/6AjwbH5dN0aQdcR7/gEANi+11Gh73xdwLtewlqFzEdCHrn4fxzutx4WSYEGgaZRnhBC
FOSt1jeaz07yWpyuLw2lraww7wK0ULcMYtlV2746LHaA3kVFp6tRqT92itFzPaJGXiM07wjFb+6J
btNJeWuNM5Hrr3oEL2XF8NAFIWgnTlIjtu3gm1QkF+yOevrx4Hz182bHTBeMN6ZFs+vaJrL/PQZx
NrXRlXiU4YF09i25G0ELqEsu+OoZLEYtsBfMyv6JgIuFki8keLDyxr7jZhvquOaavVLrQf8qPN1i
MVlHyrImI7hhGkwKSFBn2lOWi0q7/z7qpeNRI7jKVREWOzzrCrSriQgz1Z87d6wAhSNCvBPDBMBF
YRNds8mV1D5SaWGFN0RT4tJ/uXDJaMJazAHPdg8tP92ECu3EvalWj408i3f3gpQo3xfDyidTUiAG
h06gGnAeQSqTna9fqZiRW9/BHKtXLXe+3Bav60r7ZjOD3FRAL35lKvqtn5ixIqfkeTPzqakRlbuL
gAlta9Tho8oPfRBzEpLeJ1vNryS5jvWWzdk1FdJlscfQTzr2fRBoNDX/oOUqkHdTSf2BgdHondha
oM7THpBkfTDi3Tt2UA0ofxWKMx0FV8p6njq3IgJvDpN5l7X2YAcYHUa7YUgF6ccGa0Xng06DUbSH
d1cSoR4t5sQPXf7otaHBRswCvljI57inf0LdUogCcsuJ/iQdJzB2wu58asXYl9YMGVG19ZlGle5D
EfVeLzpx4mKg0eK6qXyQTJBVCQDxMrULBgSZ3fWYNcEItTQamWRU4Tzwthbi+K4ILSvAutTd2nNH
M24i+u0m1fKMeuJOzpErVY29Z0NlRAytdq0RQJA0hGpdRACb8cezK4tq0vX/cK+vcbQM7JdVIlz5
giv+yoDkQXgyeqrXF0Q8glDVleaWdreDU+vkR+V4jjnCHAlO/BXV8Awn0TGe1Q1/67HJZh/3EDwp
bRih3Rp3Ti4OmZq31idDLp1Z6z9G5UUIUBJO8sC+TexEqdlehC3/cQsB+W8Ubt6jwo+05efhOMgU
/9LirpjHx2jFMDImyJZJJykbyf5Pq57ppbUiuzyRlIwiLg+pMItlUhTEy9Gui1WneJ/eLDIyLdSO
3e7OxmRRcMewoihw/7BOLuqVDQodZk748APhALH71n94C16rwslhYYmBQuioSczZ084/VL2BV+YH
Ws8VGbUWTB9zemqnqYdB71FZiiwy5NFsl+gwOxSXDRrtPMYijs+puGG6NY4uwKtSRgE0PQGCJwEA
QF4CdWfO6myJ4YAno6qR2iK632H4GtEXFAQJ8ThnW1jgaLAaUoxJQYkHNuHqIRLzPlnIMk4+Odrd
YIYoNsb/M8rD/3mvROmzaYQC9fofTtwm2ct/x2wji+RW2/3cZxw9RvdI0y3kOwyDk/OWCMScJug4
35DIli0KofriHGbodSJevmQUbnkP8IKrECT+1CpJRnOAuWhsVvqwdW2gYMXlSdr1sN1ca8ZfNXik
zpR6UiEXDI2LUOfxIaZJK8tgJsJnK2Xm9c3pzzSRLDNG0A0gLFo/Yzt15zw2qanCdU6SihajRCi4
JddUojAiFGUFxArmKtr0C7ViBpQ1Rlk4F4dG3Zkiha1UOY0780FNZkvPCxrAKJnDFQMiR6cBT5Xb
9IrdgHVUNqzVsp8aJVaziiEZ49rvkH1Vtz35HXJc+e4fZry2wBNcSjXW3CREIGCtaPYGOm5IUtKH
P7oy5o12sF1cDqU539eGKNiXf+gZ8i7JPQTfdYUBHtiFw2uRR6Dg5GWJLnotZlZMXLWjXcxoiM46
FsT/TSsEmCsK3+/B4RX7m7wddECMI+XVSbBQD53UHlnWSlnlv74rM28utpGCkCndz43S4+bqRP1K
g/joef40bLhzbhCZdpsjTbRdAk5Oj02TYck1aQEroFs0CV7X9OXzPLiopbl3VN5n3O42+zE21WLg
LoFh3sZRz0RySu2oNgqtMPTOT2GiWb1nCwe5FN+QTVdjWoNmHu6nt6TlW/lAXYrjAgHprNeCTO5W
fAEVI2lHAth/LZQbj2PVLLsPGtc2CaamdC4T4FTSmZUOM11cSYMJF5TA3d376sNZc89gyLZzwzK+
7M0J7JiW5b5rhgL3hvjGL93BSg84gTx/Bhv8ThqdBYUHjuBN6/9gPfNLPR35G93bqPPeAFXsczBl
0m3ndUbSQw+q8QeH0nuZYqJspSdr52uK3eSevBFfQLmssXYcMDA1KRqGHvWq+9snrP+TAPtm8pHb
ctW7ZqNR/omlcwq/CT29b1oRrd9dnAtlFOTMaGIDe6qejU10QEMT5hsXFmf7jhpjZq9zD9HIBmL8
pMMFn+IAS/k/u0ZuIbXE3WxGBeMXseRyfcNOI3xnKIFo7o4RI4/FbOqIzXo8j7VbsMxHzLib8dji
O1R8PcXAqfZXYYpHMiSsgouHrNOJZTP0LgFrCosFfzK1kfMC1IhLqH9iLryVb4RQ0MLsaZYItAu+
cEd1geGfyKPsSiUolAFPcbnQRQrMTXs9si8tjQlfJz8ocMs9twwIxF8aCy4cK8FasEEoH7EUsju1
zGIB4X9scjtpZTqRgo4ex93Gn6viMRnYzjKW8psGeaLdKvInuKzYosa/9vc6mk7I8QiE5Bo31+Gl
MpaCvqDPqUIyJa96wbUnLrpmpQPHBGprYWlxAw319F8kg1BW+c9Gi9mN3kaB6t9wUbwXKMt6ebhR
oYIUvfEnd826hwLmAtH3s2/5PGX5B6lFJFTliDp49QxcuEoKfNcgZQbIUvsDlSsblVDh3BqcNQfO
2m/Luq2Joa/gHDkTpBB3OVgPmElHSWRw6SXk72G6X3G5NSAaHPhFel349tLw2dJNWiM5PRgSHCII
GxhWZXHyA/QLK/6kJcUztYavSm4IBYgoCPtHv8sMFvS4Y3YNowQpMBelfUAyn17iCmao4Bfs3pgW
j98Rv1+hlLo87QZzfXrw7eTnQ3IVxAbRIuNL7TOgVECqPNTae+CjCNKY2rJFKak5J/IpNvN0D7Gc
Ca8IbxxTry5UHih6GYjfAIiBHUcQUr2yXDj3WobwnO+8rHroIRYT8y8mboN7B9Xri9ywxEZD772T
evBkGCQ4/+1PSMGXRfTcNoP+YFI63nMmTSgIINgMZwrxx6rPIVk1HZwYbkbMlMyXMLn8f+kG3chl
Pxfuasn2zUcYo8Sg8qKJ8cgNsGhq/2cH+/K0RauKEAiXQBLnIqja7z9KcE1PejkyyTXcBWbLZnnt
8V9/gF5Lht8YxUC1CEHCKSJaE/3nlXAIiBwun0QCCI7fU5lfScOX41Fm9lsJO0it1OoY7KL6a+wQ
BLMD5gk+nyW9zNXluOcLC3DMEAcKY5mILmh5rdqT9E8DhWHvpL+fp0H5oUgMFr/8BLkJ6d1bDSn/
Jm9DrVW/ca6HNa1naSWahWL8lyzUZQ0Wm2wTe9O3Om0XINIBzl1grsaIvKiMuzNbVUHFmcFlwMWF
ua+wkCN2aj4y5EX7DeM4ksM07sEm2722aPpcSFP+wboWYPts/niVyFQnxmTxp6QtnIVx2RtkKv5g
0tGCESiCzHERXlxHTkw9QSVJkBocVRLlm6H9YZ23LRBbiLFAU7KL7hmOtIKpGrIpHYwohpt+2acZ
FXeyvD3BMFVHGvsZ/052V32AGw6aWoWpwK/PM+lrBapjOqt0Tpar2aCp5NSeX7/ew06OHqLpSegc
th1gXTlFgglNiVUjJfhxk8PlNVqr7U6uMC87AAGSUarZ2cXt6o8zf3TUa+qmaf1kbvfgtDRVwTZx
rwKg9NZiT1RFiucM6EbQcZfmBLOGeBeX69CIi6AsaQhEVQRcgsx8G0nJ9yU1F1SoaPqLVO2DjC2Z
GfoNL+IkI7HYmJesLaQTE+jKt4dab2RbBipKISVgEP41SFr9q/MK6tIJZPl7Zqnv1TslNJ4AHy97
AdrNxeW8tIT9Lm+nIyDpOBLnfcS24Y/8HPjkhfeHq52P+6sVmaKa0s6e42CGRVyy4C2ZTNhpG667
qilJdPTcI2BGSQxNo3tmaPaWB3AbGvDfBZwbsFWopQxcAbCxMihsp5uqDOfOUfPFZ36b/sc/zDP2
cxxbfdUD5Uix9dYiIojICXWf+xpvdASgyUfCRiw0p6RM6rMtNWvssLMVdajMdep9wCqDTWzemSBQ
DgF9VKQIAI4rSGvuzCBE85S2C9uqja4DvW9WMZn6TuNphaU+fzo4ig1Jc4EmXt8zpAvLouWwpo7I
UwTQZCiTQkdDPjV6rzptRYU15ipTJujLQS9cE+llbLdNOxNSahh0rcPObZtlDE3rO/qFHl6f41uU
Rj7+BG2Iy1zaAYzEF+kZ6Sjs75cMO0hjMtyRcDPmJmEH455SajnG/LuMx/SQ9zn3HIO8f33f5U1D
hM6tX4Hqi+mWzMNsVVliqRof4o09CsWqmtW6kEQN2qFBwV8byL+KJUwCupd950/s9lhCXzq8YYyS
0dYPPH+xevUlzoQsSzL4ivDRychNo3yXY105l9/B9EbLUi+dnzZrFIVpr2CwcDLY30Bcfo4hUCq8
5Euq3vT6taEr5SXqhYE4R2JOh7kAq0AbkdejYXJmemBVaxdKQajl4iF9vqfZDAvwi2OFnct/WtiI
sP3l5+cXryinhDDtnfmzST1OQZP6Yo0l+53+vCqvYZxgN9Rp0hP10BIp66PtgD+QC4tid6SJ3KU5
IIw+q0EbCbA/iHqcan1w7ytO3123R/ziY9lX9ufalyEBj/H60Oa3jQ1LfYdG1+Ruy+CZPrbJJ10M
1xEHmfxP/81qwH25ia6cPWzK/bsqs9J2r+80YtZs7PbJGc2X4n1g8lOSbn4RR7gyycdpBuX/8coC
5SIaSxrsKw1qR9kg37vpMZOewxN8xd6r+opVMlrrJdFIEFSzjVipQu0nk+hSjmwZ1JYwPTyuceMk
Na7yyJdEnYCGTO25E6Lt3ia+UwglTkoUa70qiP8HKPiKYGnNJ0+ITnaMmohrk8kvapOSjiy1USpE
KXRn52uZdREwroivsBL20mEUedQuoHIAqd9dmbFdzwm4D+Iq/dMkzTiuirRNcGFPaXyUK9UcJSFh
YCJPpJDE2wTaI92mu4El3kE0bviV+SbhA3sNKhsE+VlH9VLv3DNojzCm1pqrARHLg9ohA2+SqBt8
bnyRIabG1ZG2/blNO8uqTEIv7spwcIJan/PmcPqiwRppjcPREZC99H3cd/Jrzz8VoLWQiMU2HJeF
owpg23p+HmqCFTx58r+qiibCen2hmXehKXMXfRONu0EwaAe3RSQgmyjBuBvdBSYDN0ygMGINw9NR
s5cIEQ/DWpI6WncvDCTU54RVrY7Jgr/k5l6gkztvVPvYaKAUZJC2c7HyALZwd/beh/e8R4QXmWnq
Q58odpReInf84oVSmYQkDBmpodG6qRrTqDuuwafUieC1v9D8Am37+HOxJOxIlI5yjg8g0VTRxR2G
meKVrS7bWa8S43fQxASnhmFFYLixxuXfi++n6m918Trs6EOYe74dBTDAU3VYw0R0hAeSHYaHFPsN
DdQiNmb8BUIi2sl+tdfUlQagRNKSFVs611SGdZZvPv6L/Na2BGgMlNKfZ7DkOO07PQlQXJruu2+P
D471rMQtKqrodR9aHwL3mDeaR6VIWZGngNC68s/WFMqOj8IQqcrQTRv6XGZ1gn6owNvC8FVmoXrQ
v9/BLPcUrvyaIkiOPUe0Lv9JSWULWITJe2Y+TCsQN/rTQCO8o00WPAWL/tdF4oAQI5r2X7fv/ZRR
XzhXQAsElc/AElqCvjIhFG4SIqoBUJKesxZh0rZyBBHyMemaBoFcxf3qkAF2H6GmHpvn5F7xfHyE
Js79rg+2FATSrnsGD/PkEiqQC0Ax9qJ44MSq61abBSD+6/1TRfCMVY3C35/pLx43wu+aHUkJaWJ/
eGGs5fPfUPHjIpxq9/9UY4C9zHHzA5/cZg4tVbs4aABi6jYjAZZs8R34Pk3GnlS8EieRSql6/j8N
Db9QE7B8EdmZCMdUlo/Fnt0BeSjymxUBqDmsCyoOD03sSywZUp9KsdzPB6fQ7BYhwob0jQVXxC2+
ZtSq1OErtlvv4bDtbhHg+avy8NUvFouKMGFYEuvCuDXRgbyFKB2zKNzzBN7bNJ1lxkw6UvAWWSSQ
iW647AIJuCBvILPKtWQ09imZ6Ck0XK+EXOv6zumfuDaKjou8BcElali/TC6vWARwiUBAGfxR4pKC
EoSBlFbIgZHaBfBxRDaKtHa+mcgzdYv3CXWXon46ZwZ4RAfNY4VK7uZhVyh6aykFATkTjVbGBQtV
AfSfzqz1IFBd6Hg/yBUN2LV2wtBv9jD0uFJg4dOHs8LrCi78cmTo4wZHuxLxVqENgGWL7m14iRB2
baYNhCqThB1CHtIXJad0PttgjRvXI42wvdLOQHM7N4R7jfuF1+ryjCHbh19HExxSTEgSS44CxBC4
uzupTv2J1D85FpHLIbOq9nX4tMD53MGf1B2Y/Nul5j+fzWNB+gGQctSATTpvaFqReTHqDXbPghVa
DaaXPeeMJTtWsERkAfKtlw0RiLWIMzvIobvo+Xmq+8LIEIe7Gv+ZvBhEEU1dbE9jHEE30tLMbk0y
y0bZXxkMBzgOK48bU9wIeqlA2LgdmFM4XjAAIOmrDvOlUtP7ySrVLRfGahiMfFNXGr5K7NP7raep
v4tFuQx5RJmuwuaz5pBt/u2XOEUTMbPZDOjOgOckhn1f5JXCHmpaKbUreLWdbRN08Bk73cUx58u7
UWZwTSST367D3XxsK1ySMn5Hz9iOKTNNdjFV3z7oJwQxGvYYnytpPU0AZwryV/tIp0wNDE7abQBL
iWyjYyYoKAMXDy9ORaaq+5G/5ia3Ct3vMbI3QPMZmg+uTpjPzNnvCcuWjDBSNbb6UVzbsImFueV5
KnBLI1ywS0URQC4HVbfbKRGaNKHDOqvz5lgrh6Ym5fJxBvz7Z4Otp3pYATmxGofTzKK9Q25+BY09
UObzpIP6oaX9qGrKP2M/HcB0icRYLFB4S2Lc48IYeleYvV3kyubaVC3NiWsSwTUDZ1ck5tVefvMC
caa2jDc9iv8ykWShBSC1xy5fX306yPHW3tgQVvjgUi5dwb4ONzkgvBea22N6poxfmz1Xf90X67tD
uvVMKlfpL/cc/HSEtRfY3lZaYSkvVnXoub8naYcxhOGmncUM8YuJg7HpETocZXsE8LBuZpde/OYK
km4wMIe+hglUizsLbbjsCDVAR4A4rsMb5PAO8q9ASunWqFMFlpoj/crzPdrLsUGG/pInSvp0ENlo
ubNgk/ZZPg8JJdPO39yFzqsgMSknfPAP5cQ2lSNjN+E/x9OR7/Vvzkrit4i0HfJHHdWdA8LI3fgF
2e+jWDymAAv4L5Gv0EZOBa5ZluQ1zKgP2va9Ovt8p7E8gCZoRjNUGvOdX1UG7w+h82Ok/VJe7zXZ
uWV+5IGUkSmSm6QPThfsBPUmOAcGvn7LJvhjSDI3f9AcjcZeAejpeYrYNrVj9ZQ1aleDFUfy2tvK
udbTDly/GXRLAUKAbMQItiZU9gPaHxPix73yTGWpIQmSQkYGZmJ7tz33cxZ2qMNmt9zdkpzggYNV
NLcihtEWXtyX19otETJnz31mx8bogAm8yAOxvoeYlj6v1kmmBumQ+qV1S2ZDyKNqShDmHNrNDitT
W6qPyXMx66nvImQTOmIiUM89lFoHMFwGNCHkaMUXqfkr7kdUo+u+vhew+lMVt3jqlaTZfZlBYHkH
/HjZ0PjX9RrKxU7oGag2QMY3JetNH4zAkpz2NvV7MD9BLvR1G2i7Y1iwWmUScroxfkY7wNeEkqTA
KQtI9TKwRogFWvw7i4SusS8VoZCIjlrlaGLsnaMyYdRkYzHq6jfnR0PtPQiYOh7tVnp5vQ01LMc/
ojACWNOWH99rIo7uRv6WuVh9QMvN+YOZv9c4MUmyeMQHkpUtY657szWn0RPJd+ig12oOGqvdGC4k
eHBynb4g1fKCcGIernvxWH1KDtOOTHMHJOo7YQRgZ4l1heKybA9Btt3ZHEQW4C5Wq7UbINwADObj
9Ia/6oPC2FJvINs2GE3MOd2VkIfzrbNcE4PHUjUZLz7auaLKW39k5xWw6HA5+hSc7Z44vS7mP5s2
UwMZ9kkf658dCm3N1CE7zmjD5OIF+CIvHabrVBjaf9n7RvlCUWQ+X3EU/S3teo6mTvExNN23fFMq
Rxl/Vk/nQt09bztnf3poVMFpuaJZqMzsg1RECLY4F46mysQQOkj4LqEkgGpXQ1KdypXNgs3Fyfle
cZZbzaO/aImMRI6emhgpha1mNbhunPiW2DzWjvWz2Mx9wxJGWxXIS9oy7xHhyCbwVysTWp3vRzwo
Ao6tTq/td4QBWf0AufRlpVjGr5E+MF7hXPhykAbg0ZQ5T70QYh1qyXg6OAVClTZak5yqYypTwYDA
k67O30Km5L1j4sZ+RdaEvzkxNAZEv7xgKv2ZwBKFmKITpNQz+ZnNy/xZLjKZ5kknnmJkFcts5gO4
XVHr/QFwtcgIkx04aHwDKElhPs3U0ZccDFkSA3FDUN2JPgxpfgSftyLgi13OvthK2jt/r7HaENK6
EMUVr31sW9byRLBst2W0zsaiEpgqktgzPIJuF09E5j3vjgAOmqJjjJu0ZYhWCGFS5DJCxJll0XYc
uUO3iTYUPYezk3x4Pccu0xXacvLZ4SQZ6OQxp3vyTg9NelWZfiJ5LjwCOiVJif7DjZNyBhtMIeoz
DXGqBq2x2T3iKf90nXjtoO1Q4YgvDKL0oWH4AW9fKQPAaTVwQnrE82hwjQUpW4X+aos+ec1lE1iY
u3HGpXCfz6wvmnCWWk6SJhTj5YpfVgEmbEVJL26s2AEKTL2jNwmnNGkhEByzIXCrTz+0hn6lTss6
z//4rF+Z0eFvUGDnxZAR5+Gq0qENopZ0tKgB2qHdwWkepOPPcquccof8nP5WYMhryf9Cm1I7aH2B
+haU+XkfJfpmV7N3l50CGq/VM7numiwOKAsFpYk7IVSApxDymeg0BSqiZZPVRue2PaJS6IZF+03X
7ZwjBrYBt1zckdkaZqKajhKlvhVTnbf2g2TmZ5kMlbeDIUaRrR9eN3zbXX3Mu2D5N4z2+ADu6vwj
wh36wQ4QWJ1Xgv3nzQDI2MT8EgW7QIrtp32OBIegdzP+poWhIt8uxWy6TjAOvcENcBSvZSbYIybz
iz8eHwNXxxGYO/MqwxiqkrAjr9EIRJD3BLQyaVt6YZxmmuBpTapE0y0CBy/g3bPfZZEuE5wZ4fh5
gBmemUDufULrLGGpqW1ZtvogJ3h7U2iEtxmSEcfaWqGy5mO7UOo9s2vMw9ncQub/EZo4oGzSHxxV
kL90T6XZbFRSg0mkEQ1Qrp3H213OI3C2Wh69QO29/WHT9jkRex8uZepC3ffa4CUkvjbR/HkGIg2D
Eb7Tp95tBhUixXDxX5mTvohHzmgTKYIzdHXpNvaNyViJ3hEyp8xHiPIWBV8n0z3Pv6nXAN55bJ5G
95t8IaVeB0rwpFZumh3zlNUKXFS/y89h51aJBnyzl5KT7KMwhFwL4zq3Aj4LyNiArz2hZHt1zbqe
rVEjBr+Qjm2LsocrPIFLJbl0U+jzAdnXZ1bwVUPjtLDnXISV1ScU1BGvsQqiJkx4ml7ZEcMza7E3
smraOOokPGynMVAGH43bcmzKS4ZXVMvDO0Va3IMy66qaSXKvKqAR2llPXYWSDDvukvwk/7gDVIK9
c/x+58whUpb4XP72k+eJ2Zq/4j4zpAqybJG41k2oCYYv7PWSOrMwZTuC1YDB/XMgG6UXn2owe4li
GHt+ttD3CvLUm3jCOH9AlEW20aVb26LDeQ3RGLFZLjs99xHqdRgoS5u8nnFIkdKDThXPZrq/dCd7
l7+DB3VnZ7keEon3DRVrhqBxI5wICIthQE5SI6TYaoYzjJR2+996qzgPcoFyAn0g9SYRgpQ0ZEVC
VlGtcZIQh/PphPKfCcumkJFsjUFRdDYhyXw2d3hZLp7zAoQa1v5u32JgpvZ2B3IYmFiOC/ApKo0u
+8obPNsQVYIuN9oEjqbB3kbpgTzwosfyIQgK2TcRyX6718xfqez69VejAockwviHIYhK0StcFGce
Cm7fZwTyWvDKurUjvdgAs5may2vSe11HpUxq9fTFR+OcNIJA+G1AXn2FX2BIvMAYi6AAO21wll8V
yncY3XCGwH3u84T8vFqcKxrvEZMK0XN1P5ufSUoNclGMabzQpR8WwUScr01UE3cIM8dURXNIDO95
k+pjeBfaEgYvUjUX1oJOebM/wuEhMAEFCdceyd1Z8DYKHjj5Za6WyeC6twOn+ZUt5sAiYAtMjhTP
9tPTvYTfI6CLnI1HyaOcdgzobQK0v6K3UEAftsxKYZhcg2pZkaHlFZaBUFjRBXeislfg4Wg9zikv
+96g88kHBjCoBg0E/KDehnVp79y1F41MLrjqAOfqiNOEjaI0ySwOrdXxoyAc7mzulhIoayR9E5pq
Kf0B4iwal04kaS9ZixImCCtyj8S0FMmEaK2g6EgAHEGksaQaDqbuYEhTRrNlEA5dqykfrz4+8Fve
dtoCKQWW8tx7iWOsfxYY+JhU6GshK+AiendWGbyDXVy28LDL6MFSKzMKEdyE71M5hY8u02KC0jta
DWRil3UbVjMI+h4cyzOaUFlXPKXwFfUWIEdXDM533VUGSfkqZQgAhdvNbSfe8rPUYPXh6yyDuBWN
LaBHiuzBYxzWKIhDvXqszJrnkzusMH4cv+iZKvUidTmmnBopQ8LGeI10v+PNTXsRe6G+n8K/P3nl
Flc7/3bLsUqou5BJbfCF6fN/22LovF0MHTfMxeHFWfwvID/b/jsdIzY2u2LCyAGTwAvxCEbgduvx
AZvCH5wC/T0qik0S9Uw1V02G0PFUOOxYPTYK+Wq2aBpCrwDZy36Evzl9PIpfDSbQuBSmdntCkLNY
ZGa2sn6d9dj+jqSjHA4fZ6pVpvNTGsZnU1ceUztE4U7cGpxGLeWSI7hfNhkuDRO0Zen2umwBxCca
Q10wmCJJOBk1FAzcoSsQ+v1jtkNzoiDALC+bRPAnkh+sIbpMOkyBIF0BQcffvkQLIcy3FqxtMVus
MeYp6bY90ucUhKRk+zJP771BpGg8VcvO0WxnFwtNpmtFUOU5zgYvVmpljhH6QT/zzwtn6H574V+s
GA0Nx/A6nMU/XMdcjNI+3mv2Nolfd/JLWEIZTjw8XY4bCTrXyFcUsJJtN/r6eQZGQuDLU6P22+F7
lqXGPbZZBN0BydEIZXOb3z1/qLkfFRsKsbCQjwN1ToEr9XvQhRFDB00DAqoR/zhCsJIc230UonnU
VWggVrKMCZ4B/wErEkNQ2PcZQFlLwQVTnmr/rqAMaFRc3T834mTu97yO5vJEIS1uHr3CK6UupMNf
mJbLaJGeDL8cGp0iHKBmYSBXwphPSurVwE5uOvt1y0PslTgbjeA47Ci2FyszsZDIJdTYPFM+r+9F
Z46MI9en6gdChCuF1qctpgX1E6gc4NW2T26qWD9fYHG0JXbD5+dNIlMwvTLebj8fpU/0hj7NgRXA
B/cdPEZsi80FMdjhSZgcekK7szjAn7oO6szJjeZblgMd63xTXxfQWb+UdJ24VhfgU9g4c9CyWhN8
lMyFsEvMb+dxd2wo83GoE7PnGhhDC7FuwY1IbuQ5o4Rvzjj8AoKexA+kQRSbVf+v3UEf0URSzUzk
D8YrNM3y6nvYJ51MmMqlhUxWAnl6fQU2Nrq8FVaumT4cxR0StPqSIjnw3Ym9kqlzcwey6qmoMoln
/ImWcCSnaS9Kks6nSCGFq8EAdbhs9GakvDqIX5hcWCeGnBcrusX7DZHPv57TiGdJhdCoI9WNop7n
2jZNRyimoQUEktkpRgx4IyrAYJ7N50d2G+aM5RuqNNjSuK8bFLNfP3xWtlb3wiuUaa0warVMHoE+
65LL8piK6Odd4AAD3cXqg5MxqzulT/8BllBYa0k4mxMz/le1Joc1F/jcAOplV2IYiR4rYwGxVFtR
9vhtwOVmNuvUdE7bi3TXTS6pKlHzaVvr+e/2tGIn8H0f9a2nfQI/y1ihqiSNb2jO2K4SvbCCrJRA
QoK9l94Um2Ayhum16sU5EoBILmPgiT+m0j2fatJofJjBAFcxHKu7HfuDOJSvD2CXzvwJTYtQg3O/
64TGltPGrQH6ahHVPlqHhxBXa6m7K1kYTa7hHsD3CqIUOvUwWSfM51klA9TgOadQmfo81gTU1aAn
0y+rpez0pcE+2dCsB6YNAK6+VefhrivYmDyQZjt6k7vSg984Iq4fVLM0kZckiB/f9Vs1/WuR7AKF
zXmK9LMb6Sd9I6bSYVxUPh6oRXzTKiP5aaJwZ/5OqTry9dMvjEhqilpb1xlG2pNmX8YJycT5N/sy
pRiiK8zX/ig8aBJrOvRhpB+/xd/mRgWoOwcD9ZH+R7VDEoCvcWd/o2IY2lMmDgZypNlwiKMlrsd6
sBWdYdo5TbmJVH8120lfQq+t98829BhlL/tr7aNnoS30dsK0uMNBcGcKc0gd51a+5NptKEt2H1uR
OPA3bFEDTseFevPBrQSgCrdkM7TPyyCRZLYwW+7R0cvPK7h6+X19rrwWOXjzgPC02XCz1KQaNo7L
/Z4/INDQDgCTXelaAIe/dNCRoqLzkBjHVlRiMsthR/0fY1L3lMBklZMZborbGvEN9EKusOgEv8zH
bKoajHTTl7+e1Cii/DHxJzkP42mPUqMFaVtHRiig+KuJWp0Wh/zE9zJz3nj41R/DawQSnIhY0n04
YU3/uVBpQpu4EJhzH47/2NoMc6SPWP5XOpntRkfdHVBWXGQPdNH8jisQ03yWJaKgDAhXZYBlIp/u
lgzJBg7IxmjL4l7LYT8xl2HmuI7/1INAZhIH74Rq0bS5ELvw1CgSBabRYhViAiyb+Y1VwWC8Sxeh
86Nh0onqhsyNH1n25aMwq3IV9OFAfxAaEyhgewBR3TYwjkQTBUBzLAfatkqxfN1m829vGuektdTz
vxpBQLW0DfiBnfg/DNoJU6Pgymq3P06chrTLObrjDg5mlh5bmMEPiitEp4VTYZC5G9wFx6axuOBJ
g2CoKSWFJAvvURZK3Vff/J4uWYnNf9BEmCHZKsGn65LSJyoTHji4MS9b2n9CrBgHihvVgFBqecQw
VKcJdkPFuEymr3RVT0xpHDG0nmQbijEUIgrajKFIziKrjjww4GRO4Wsh7nMszaCrM1GxaHdjTKe2
XaWcKPon0c+brPE0L6mAmLhWOpRbF0LY31jzT3AX9gK9g6MGoufLu1U5WAbSO14XYVIP9Xbvk5xb
6zQ28EiVwu4KsXO6XMjunFhK/1Q8NFDASFW98o639vXZGQSWHqQIdLMk3Xc5kvJR6Trj9GWkZXCx
BWivNV/nUfth0RiVrzfrVMJexID7PT89KBNeLVOWZqC4zxN/5mp20U3bKJi+EQ7gDsO2w9RiDDTk
TaBF3b6Gufz4z9JQ3S6m8LWXAMo26KJ27nfXfmGNvCUc74YBNze7vb2aQJ61LoVnrgxgvbXsRRv8
x00pD7N5oStx3l83iZ+zUd8xI/D4YgSJsXnBqR0PGYbfFwtSddL3cRBTS6I7lw263wN0zctm8mZ/
Uq2vW1i+iX8jc7FkEoBiQ8d+wGzfICRtAM/8OSfNfWh2056hwfOe0DB1h1ztfkwpDZoj4dgvxLWz
Fg8Kvib2VZWIqSYQnKMcg3LFiHBmF6gwliNIHqdWiWcXAbLZ5ovVnI5T7x/YwBMtmN8PujZ4yCDi
ur3gohQjq61KFSwJSHQeUmz2OtL8o0T2U2mxo40j/96hwgmRdIqAi+egyzx8heK7zVTl1caGFYcZ
35b9oCuS1mRLbYmfcHdcAN/OXSqZrxPegtcHtxvGDDxgcOaYmitmhakWmZbWvaQLpDP+4OTRgAZ2
SkRQevGXe+8tPxzh5xN9K4falMLQSz76uSPs/BBGZF9lWrFf0LyTO0nr+o9wZ75ZIC8ZvcBe3+qQ
vHesvd5FboCHYjj3P/j4pDib7+G5fQSEIHZ4Ijbo8FZDpFfDDEyg0Nlm7NSIpOugG+Lgw0Q9CtAF
4gL695uQWI2K+CZjk3yErees8YrvjpIRQh/IYn5sY8QCiHaOO3e6cSeqjDeQTAVH3m9HZ/dThFVm
VTZMl/Y53pGmPAC9Sbw03Ae01zwUq5OkykXLh1r4vxXjMQYzt5aJkzZX0Ccd87ggaj0J6JHtNGi2
GmN7YTHBHI1pRE5jPxHJk/sM+5uf2/MtGJymKoDdjpMt4A26jOCyZYvXYJTx7ahgyHIJgYPWi42B
6wKAWMuHMAwjV7/yzbk4Ad6PeGci3MnFme3a1xIVIftGJFseQjWloTn6SUo7IwNTPsK3Ag3g6iZs
0+EnSUwnzTkKvsx71FJ6rURx2Qx3DSwP3t0J23hY49r9TieLNZmkw+dlzEYAnhuqRonhiZd28JHJ
J0mgZsyWU2nCr2qqNZtqJ5EUEB6U8zPG1bLxhi3UNs75Ev6J/ttje6tTS4r1HRfQJNr2rriFMZ4m
qkLG4fDwDNekortmovTnTQNZLw7Qzxmy8vxHMxAdDQo45XPaSWz+mbNKtvs2qf9HbTa1DBLBcoa1
PkBr3R9s+XTg+4ZwlBfNiyYFQ8NtRYeMEMpy/bCQ4srYbhaD5s4o0DoUNgbk0ovAdiehxVyA9YIk
/9NNn9T0z1Jdy/lLte6JSJtgnZa5fsxmltVYxbdBxuS7f6wkyQCY+jJfPLVI71t+sCYHujb53DHz
ermkibVtdtJWYV1j8KTrGg2aKyZtg45/dDElIZUYD+fVKPNA+XrbD9ysD+RmEWGjbGuqMn8MSQW0
daafTvk26pSRu6bAdrW/sFA7/K7ARyor1t4sUnlvuKsD4Od+1Wt84UqYm099fgH8wP/4ALi9sfIX
T4fujALc1tAAn9sAKM6nT5Ono9Ru7N3o47YGZcjUpO/Ymi+IQR24qfIEL4HeLNgCm2dRCZWTZYSE
2etLK6C1j2XsEGxxhkBeBYz4IyXnfBGJf0YSfiy8mLKI2/xn686e+WszFdkGtUJlGS06RWvdgq4j
Ysca0XbI4oaJZr6+8ABRLryS8onKkyfVFvUuK4PkkZmedeOz9PODbLKtAh3Iyot/Obm6OJZjbj28
wQy6Dovk3w7FVkJPd87Uyz34gGka7hBI8zv94nbql2gRu0j8fdfF1Q7gzA+EbwLiVrfnBctuYVPx
k6ZK8esbnbh8QsxITYyk44U7BUIcMzbWcavr21CVCH8ZhXA4OXYrHNsHjVRZTg81yRUCU8Ckh7xJ
c1kKB5u0YA4r/CxPDnphEffLo0WgtPHM0CE6cJzFgGuMLCuC36BXt+b5ANeWU85xzPGAanzbo8cg
boKa2hp3e6Dg5GtsUU8BzD9Y2gH/pBiEVydZCH7b6LTqrUYCeFBen2BzJAMaqFzMffKMMc4+kQEg
XfKgbVS3485ppq5jv8SzVh5zdE6ATK3VyLLSrHrVapBwKkOyNLdEOUEgYHad2j1Qw/kEpt15FD4F
i6aiEOBjMOyL/c4L0ODK93+wM2h0aUqwL0vPQZrg2Z+mHn3G96p/MalGfkiCqk6wlBtg6hi97Zoa
fKXh7AV6DDn2n8LPNCElkOD+921O3/nUxYZdfZr5jdQ7Cl6KGW2F43LDAUVkPovXo6deHbuoFsTr
QYu4w0cqj6glf9G90sCmgrqtFRhxAYkGSrgLRLE3A6tx7AiXCzyCkD1ry7PpoBXTjVSe1yYEKM7t
77wYDFhALANrHl23dJDhmZScOZXYR/NYqPFOnsaqFgggDUae14sHMwvLRXQY/UlfXmRVkdgbZHKN
QRQhTBa7JCkl+rou5DB7dz+PvmkSN2mmJMEKecvAokp9duU+Q033rFP+lhjY/hjjdLZc3GvzhOzZ
NGdwtB+OnhFYHlhlB7iGepPB6eD2UEPWkVjNMat2A/lVx7g1NRExnmLTNvZdcbtItwutvl+S5E6F
E4Ggof9k+nJQ6sXRGSMT+IRutSrs1O836DCvrz9KqI0Bufd7OZ54RQj+TX54CT6k2Il3v1G5n9ht
a4RwqTI/vGXZ582Qbt+Sv7r6/+nkmP9PgmSdoiKQb9vsOKFoi0+rsetEokg2Uiyqo1qLSKzzA/2R
ZF2Y49te8ect2Rdj5B1PWGsby9N8GySNIIhVngdI/lxYd2fw7/C6PZcAspUfivvApSvwX68Pzolg
1FCXYjWYoA+QXCpAHviSnxgIi2EMRTxo+yg8do+QzFGw8zK5Sit83AgMS5fCp86+5erLilmPyHix
M3cG5L3ohARg0pCGNuib5anumYzICH5sVuvhNZCbQnBjTt86XFgs7XzcrA4egDCGzaqq3RIlf1QR
qGI6iyWosd0LK23wuvKhnxCgZlU7PdhQt1PMGPKX3V81dZiXchhjX8PHeFdOh5Z09cpz/zJqkeBc
KN2NVDcGXZxCiuymyHh4J+DM5kxBC5F8pvNjt4RXb4bpIGR88SQb9Du31WmEaw47olmdoppVhs6l
FDJ4hpOB6UdRN9DPdnF03ePulpJmtGpt10LiP0hHT4gjSsBXyktPL8KeZ+EmpD0y+6/3EKEk46JG
Rre5v27tLOruVCAi3OTdEv0Ef0+aldko6+C9rBzDePysj7ECkA/lslftXwf/3f6eYkzh8FGboTK7
wO/i+AL0TczWXhwXl4MbtRjodUoHfNv6JtmNyLda0agiIeAyNIj3uHaf1Hbe0ocxMxEF7Vwgc9Xf
YqbrYMDFt1RPuMhkVfl34kkBsoDrlB2y3d9ltJ/ul6bdFp2xLjU9KrICI0OnRr+3Ifb177pD1Fpg
/7RxQy7Xe/4oOOZgvh/5ZlrmH04D+kKLELZMV3Ne7e5Oh1BeE74D5N8C9Azeqf2FEDQWVziURjSt
XWcfSkzcIRJh+fcIPBVM3QxnPdy8nTfv3hYnPvTaIge1wXuUCO4kORFsrGcvqmiRasWDXmI72afc
TGWN4pIZnLk800Z8PCyDgEQXCtXSUfxy8UXjor0cyLVrkRhIuBS5TSnfT9ob+iU80eEWREV2ifiK
3tUEv7+/pQYHkbpEqyhnBGv1CyfRWU9vRb9BJjUj/7rwjrqLQfquBqWTtNWZ1jwi8GzBoRv1tyLJ
ggRZTO/Glwucutmfjr/wIyuiIL7kDlZ4GeTrz8RxySJG5/5crBpgZJw/Nt/kUvDNSxXtwgOAojJL
mwE6I3EtBi1/eOgu/HE42PMXgiFnSSJqP/EVoo4EOudYmOn6tw/WPSGl82O8M83wuNXOGlmEVf/E
Etg/aGjPe+/JwC+DGm1+S/Vadar6gsqxiI7VfuAN9sBErnh+Lr+01459c4780IaY9/EOiwwz/utw
tMz9ZpbMj5p9j3KMAzMJKWpZZaCZnS56KyZc01EfN6FkED+6dW/oxUKWeVN2w9WRK1qGa8L4E+QG
Qs8c7yf4Yad8p4JZbWKvVmptqCHNP9/KlKMfrbdtDWhks0oFv2+1fYgNtiFM9MNgZVNe3w1/cmJw
tp/xuuQ5rtLj79DIazFj2Fn8N/A34RiE9Vy/eYiC7JmlUC4t5WrwXLTnx9eplUFJN2DZMXTTjQKR
26/0W2CSmqA+VEjftQzKgcIDld6fazSuNDihPd6GCyM8Z5QGPce+XO/PL+5tkDpYYayNlr3rZ8T/
RagDhXe36Xccb2d7Lb6Ci+v8aghrq9GKnIQbK319fblmsIxSwngLmlwh4imm2/VQFU4lNyzcvYUC
kM/dkEoTKb4mZSUFKDUSnUCenVpayoayXs7mWI+MSrFPRniQJ/jEG82BqJ8IrIdAGkVh+fL8O0hi
hz1PeY+qIxbn/JP3m7nH1jlLUM5sx37HoMiPa1McIroSqXf5Hwfpjjg7Zyel6BGaZZTQZcShzK2K
Ohfs6NB9swd0iVS/hiWjsUok/7sTU9t6kz1RyMB7ltqJMyB1YtcUp4eJLbnuIhkzQienJ4bkbIns
AyrF6ep3MVy2f0keX1o7eMywlKYXNMoKv8g/jo0h36KxQ/WmuNRer8H+OW/Ts0rc1dJ55IVnaOy5
n4a6ls/lY2LW7dlSZ1Ff59MhSe0ATaI90WGA2FO/LqFpMhFCrwjh6w9OiWF9lS3EitbAnivx3aja
R/CSge+D4LBdNH64c54vxwl8yUBaL0/f687q6EzZWOLddahBoeoGgPmD2hjqF6U4MXxZ8oITb2mK
AeK5ZKtXlXMuHHsvmxT3HHObSI5RaZm+2oKvRQEb7MsaPlHr3+6OUKlZcb30JqsiDI3UhSXYflfi
Sq3F2/cNEC3c72BEd6zaysO+VgANUaFx2swQzcSI47d+Tf4RN8Mf0R7LzkeX/yr9nueYdao4Y3Qi
X8CfiWHerke9R1vh3J45+JQdPu4JfyJwaPDbsfDMUjM4J6r9AYXhmPCOzVPhNewliv15jgaeVTPA
KefVQ55ULuRyaOp2mlgrz0MVLul3YlpYHsQ3m/OxkNcVDGQVSCPeHSLG6wqlyrDfybGPooeXzpqH
Hv8GnmaF2xC8O+us9Udp7bw2xwdlcGIhoUIYFCZ9JFT8hyKR34lvzpiRZ9AWJQnlPgLqpxvh/t6y
thitq73o05nVChQHduZkIYPQWfiys1RqUa2bd0HVqfBzW5ER/JqWKAsUaK/oyv/XfIdp+ThsNNDT
xYj+X2QHV4erDW3YmUft1cqpPmPCyPohyrrpM0nW5HVMZdcT49oSI+e2CNyut2FH4F62/MGaLTXX
pG4MifdBnV2J7annwpP9PYo+t/bnXsASTUFSYdBJAE0EY/R0AbvucgLybnbvIRRHdBo/Xe1N0h/T
DLbGHa61awlSIKlV9glMTbnSgFptmDp46NGPfQf20Lf1udSue7HifCjIlNDMjbJhMw5w8t+3ls/w
G0/Jib4HpsOiqhFv4NeHmf637GrRk+912U7BZqV4Z0txBI5LJqfqyrIEs9wiNvBSjGpJGlMPgvIv
dGJFzc/704kz0elHCbcjSH3OM6L1Bh4CsobwFHZyxdgdgKTgitBIBGGx1GRjL7En1jtqMmpGrfJ8
SbZ30lk3Q4f0WXIAYTt8sKzXnkfDg01rFVf02Z3Sjmlhlq6v47cakjIKMWRPKqYLRI2NzPRqwqvA
RsnvRiQAX+oFnSBp6vwrutVdU1UcgxRTCcnODjLzIUAy8eiNUjpK6Zmr/PieeYDz/RchJuJPXDVZ
f1Kg+d/7uBxSjrI/e4A6a+b/XFosL/FGXG7EfKmvrs5wbLSzMcYxLmw2eNVF7vSsjC599HG0Xpep
vGwfp75DeX5ben9isW5ifiYHF6z6HU0out2HBWI+4NFDiWuQqMG8K30ikttaHdp/Ry2nkioWsR0P
wu0o0LVLLFxprQligRGfe68W+hoQR+mQYyqR70EAodzydkW4NOqDUPTwNRpqFzoapv5y9mLh1MMI
uPNLeS4Y9x3szwFVLoR4l2kd/Ym7IhUsnc8+0YcSst0UVQcuWWe1so9Q9LheFM1xXNfG4JM+hrij
U1+fDbaswZr3b9Oms43LelTKRIhyFoAtA1E3DkKqSRYXjYNie8O9B1CUB/9B3IapPfdLppvgTXNh
6uLIxub/q3DONYGx3jPJE4/4tPGm/LTLj++Wfy04W+TlqTLujooPjzcwNFpZjUdGRCmqIQFFEiYo
XhO+is9pElqdG4C7jcGZXzM1v7B7Cb7zs8dmyiGy+leDNO0ff2Z8JXAnB8WlWnDDrpz3NIvpI52K
6fxM+bk2utWgyQBD6UKRxePjkK2Sm6OTaqPu9+1sp4Y3M6msZHfiGE0Mb93HW/+a4Zly80X3CVG5
EhE+b2SZD8LRzHg5vmt3B+hyyb5pP2vsgCmPpHheiDygEPFW/oh0DBAxNTEMgRIhlg2qeMFCi2Nt
fxfnp3sW+70mmn+7ulPZ0mtH3Krs2HGPG1EqTd4Sa+JQyv0CT5pc78dKfdVDs4feMwOmNjHVuJng
oT/K93Ut0ZXPfO0EZzTyNzMsdbt9meaZnAlEGFndIEWhESINLkJs1uly7b1WAtTbSS3z+3jMyHmy
Zg7kvegKi8XKoKzBKZKzhrC46nju9X35ribhsiCuorW4ucEZiTGd6qXHgt9749gsNszn/4kRuzdH
QcxTNxsz5Xm81iCrwOvHHg1u72JsKgYH+ljWi5nSQZFxG/Gt9CINQMqxeHV7WHBghTyjmYytIQcC
FeABCX/24TZz+XR+aKhwXHheEMSKzZN7Nn7T0oT/Uccwphfrm5pfW2kmhVC9B3jtVfUU13vlx0vR
Hd7LxvXHFfvgMku1t3pKmulj4gZGnsRtaJNW2TaUe8IJiRM/lekTYPQNKalGQQcCD5qlHpnL4san
UrVmzuEugzjS6X+T7LmIU4myAbbY6txpvrtUF6AqVxempWeN9eTBF2rtAtuz7TyNFH0kS6d4klfm
W92iqxwn6bvEY7EwMX4TEzaPnFBLsmD0ihNAV2N7ImuQPpiN1+zAgjuVo9Lup4QsAPO2ZxffWFzA
uMMCNXV086d7sRTCJbgjMUunnePJpjo0duiL4bPpt1Ka4eq88W8oiTPHnagtzDZK3JKBF3+dIXLC
9a94hNJpFDVq6DwqUX74eko9HOSmhcLtpxe/UebDPnqVZ5/MdapY4dINWxn2yHaBd98R4E6DQkMN
QUgo7atiezSDydkwxOMwoqHdCwr8rZ/+CbDVesiP6TH1G3QoxIkGsYivKKb5tXeALqDo6JYOCtx2
v/QbFWipQOIqzqxIgJ+elfQUhZmO/u01JImmuQj9ZZPXrt6ObAxfTeIcHkBvJ5EXX4j3gD420YPl
PiZOSw59F0B1EyIjfRJMSeFaFGE5+MubhbfIxetOvfGp//CYjv97wsSrZPTh6ncgdKB/A24o6z6K
0WPjIK77cJClxGp/VqAtiZGSUVnDOXcpvp19RdRRjif7LKDxN6XI5dxKlRX/wlFjhLTRhRB/Cf+b
41W42hX6dsPC3gWm6GvfNPSNwFkM3ehhtGhnsFvS/UYXFKtUmf3IMHmIBCf7vkkS9P13G246U9NR
4JH8b1GDnL4948PP079wuCqBHBcM1rcrvTdu2ujjeqjHzryE7q43arpRPV1TkWTNsSg7qM7gUZ6L
jIRE5EXQNgYTcfK9RRQbjeAvuRfxHKnVk3ERP1jx+u5Zf5j4ITKn9+ShRTlC6/JXjlEg46y2sa8+
tScZwPkQ/0YXNiQ3Gsm1uGJFrQZ8Im4BqodkXwa8eK4DYSo678BRPo1KfV5gW194YKW3vz1ug6u9
S+Fx5uN9jERYPFonNVG7ZlvtT8TJ5nl1MyzTEM1M/2FwnfSwO7cWh8bb1NzbEscakWCHaAk7MDEo
L4OtRY3oqy1krYARFhGOo7rCz4qaUzOcEtnNimR1lGpcM+HJTJZk++F0We9GsAY6m0jE8ORvINnE
AqpzzLDfM1LyC3oQaHhv2QEvkw1IN9ggmajAsyIVE/I6veX5u9z9I/RTISg8xc7quC00xXUl6pA1
1AEUgs98r6TwokG/Z25lDxE0HwOavutSVOv8M+0hQ7/SxTailjJIORgkauBQ0TY983yL92GjC0UH
Jg1c9y+MHyUhXGn5CJZmJ8AWFdbAhQ3+Kcd82ZK8T+bW/3J4Nv5GEeW+ag/u361dFsDh8Z7uy9EJ
R+1YKBs6nqEWSB7MqXuo0IE2lCwMphi+/jO9QvOHfqJx/HUg0wABGJdvpMmoy4YgaU2TswdFjigh
CMtVGkkeeRlbgc5OWmZSN/PksizHyjOmhxfEoMndXeiwU7lkgxVupGE6HRq8hwdyGei8D/503Lfa
SW9OyY4Fuk+s75n3PghPhx3TwG5AsuikWB0Nfj+pOUBm7MMWQ+G4x4TqReMou3FTa/lvz7DRh/E/
tUavaXYO+XBiGDHCHjnj8WILFayUjb9Yc2gUZLCSxXWWAyxBBYttszBpuEVVV2mMqAh2TIS4CgX6
i8kIKK4CHxUN6SsBgWypu9he2K1ZpqolVGPElViKUfWBbey5AK2TtlvyZci0vmqzm6572GHGFDa1
EDPbw2HpzmYyS3u6sMY4EEsZcMclYn/yrIAeq94jDaFVqa6RxAvFPrCDTZPZTfneZZkhU2PMG+XT
oKjEvPpI7j3ya7Y8kn9oCDKgxyBqYJnKcshCnlaGSvF0zfh0UGe96bZ+UinCVqbeYfoc+/WslF2Q
MR83kzS9dn5rO/FhAl+r78KMDqixJSQ3+AxusDLDhqDB5upEv7OlrV1eeKkWgv+UKZF/22YbsAty
97gOX2iWpiSTWSbFdoib0O1CI35of4ooUjsg0PgH2ayssctkzzhzkbr8+mC7SFyJsPCiM25T9zo0
Q79W1OWmP+l7mNY4TutYDehPg9LeIIri/hUxVk/Wr3nFWuITxb5JHHh1MigA4kmB++YyvYXZ4ZeJ
wGi1Uc9tZMGwMo8KgBQOu0upW0HTjhx8YaxjigiKKnEXMjtcVf/Ck6xfcbz+LP1Z8WkTvL7+RX/r
9tYrzioP+/yMB87CWNkI0fBG1yt3Jubfo0djNsxlfVsBAtDDgW8ANEwEkqjMaAVkNtffuWqhy/0h
QVP73etTee3i/szGwwfpGYXjy6Zh5FjkneUBVvYrjpFe1IQUoQCfY10h8zLQBWVKk0g7YbOl1KfW
TO5tqFSoCXhILgYE/j7ccE+wiAnmUKI5s8EkkgO5Z0n1EqiH2EldbWvjx1o0k9S7HI+MoBZBj1T2
h2t+YE5ZfbnPsBxg6NKawTIUJP65lONr4HhFEngrnlJkIsN7ZpzxhZc/LZZ9gVQcvg7mJQDVyCZi
QkVt+wmGZp/w39qzpuZ79K+MNh0g4tvpnOzBw3/F3sZj7tswG50k4sBkO6rCuOSVkbO/UpNLdd0w
iYCgO9CM7AMh59/vEtuFoTM/1r8NEsdV/NqNS9DVt6Ed7qmALNlovpuYi1gU354euqDI+PMk4fc2
kvnNFOk0+dxmGIh0AZcVjvKn1sfBoAZ6JYt9yEkW0I4fzF1GFDMFeI+EBVpvbyMS2Ya4whDhxeCO
FaMe0NQ9f+7zyM1LoiaepGvuTUj4AbMUoCNrdQygif6DrDsRbUByw6qKaa3xtUTYjhCDjn9+Rk58
vCgnEMSFo+gn0mu/ovxygyt6aNYTsAdjaAr8+U9+KtrQNY8YRWF7T0guZSmb5s7GCNmqMtkIu22F
Izx6jHA5J8YNCO2WZ3mHCTnuTNxO5VVTgREjtmXSMNqAJBzvy12V4ZGuUTYBGnyZkXKeNDzPEn9k
SNjgCmfGN+a3sFdP5/1fPWcz6E+BdlsrlOqCmO+a2KCtbh/ElaP9LEbkCG5wv9pNjUpf8pgM23fD
N1YJbfgCY6lQciWSqtehMEwQ3rq7NtiDtsqpCKlUGuyMKt/wr4J4m9nY9n42gGu8K9InKePdQ/2n
6ifNNFcIiZTdGvWnwLb9essu/wjeUrQuDttNHkV7x8yVh1C6MMvXRR/I6+PhiNw7WT0DdbWENGPy
kjJCy1QQFdAtIIcJ+Zrbc4z4s+GCgHbsz49SfgoWmQFSV6/VZIZ5NiB5lyl7f2TdolESI2jhgXzw
Q5WFiKoFWtveARJlVUPoVGMZWBxPs87w/H4PMPB37mh+BEuq1aZwDb9+W5htXZjrtpkKC6NUi+Mh
yOS1zK8oFbvKgMaVR0bUL1sTn5dmF/pyN9KFqYGMzMU7xDJE5JrY3E4vpV0WfvoQWEbIZTBLVk9C
wj6C+Stsna1og/dFeFTSmBr1q2pqisR4AsqSIOqMEXrE3a61ZZBibiDRdlftz4SPR1OhrFuVve4t
wkSvfcWCpZpto7T/vObO0Qqc7FvcdPxVv6AM//GSecdo2VWHmkcpP3e6xLwspoGVZ5HUZVxgO7Zl
w42PWAtzP+U4TqeCeVWbFbqRpdnabZf/hYPGCdd3hB3O69n5ZorikrK9ntK0SqwuG4GqmZjnOPxo
JIK3QR1E/Cl648uljmlHUCKaBpeyJ1D330cHy5vw5yPmLxwh9QgJ+zsHbzf83jO6QMXgYIycZjfu
oyU99A0gzOaGPjeHJ7180L6zOGaC25GLQH7wWk8M7hct9n4yi0r+YfXnTMEibrh3oaz3FHLRnLLK
xe8tvJ/Tt0gMxhEMOHHAQNAUXijlEXDVY25GP/1f18/Z27hKaQ0VG8CTnCP7s6LgMp6o0MRNXi7o
q7coZlmji4r70r0KdXBAQu8LiMCumzCUPhGQC4jkkrHhj6hl0/R20S3EA04j4J1A12nUHnLP7QyL
t1WwrXChMYjCphPu5hgRGPPJVaokaGEhjTblHZYj9QfSA+PS+CynEzYUqxWefLzibjO98RNhWQt7
W1PAQ9XNfuZwyI900geM6LkgUYVaLDRzlScAnTtoVSKU9aHiwchjyxov6pt4atu8DTBYHCaOA1x1
Bn7/hR0L1wSf6x81DETJ78PW/21s53azEuzedRLjx6JPUCMKxQtcbVPRDP7yOKdtdTf5x9NP1yY+
YXqstyqUcGz5PhOpVc8xO0jRIQOgJJufMfjAkelr6/CH0+rg9OZBTlNLoZmp3zusc853Kn/3A55B
95VfqJqcZBJxmpXEhGuF+cPivymnQHKeteuUwIJ+EatPTB6sSuaFad5Bgylwb0we78tdR764/dKa
uBVJHuuz4F5cF9PD0fs2mFY33DZg9QFE6Oi8haKOhxxhqcrU917mzn8BdTCSk6tXIQHS8XpDx5gQ
seKe9AYZB4RIOdDRzdQCPwg33Hl8Lp6FMVkq/dbi5BEooQUzLyk+s8O5Q2McRkXRrUOMotP7edPE
yaRV/WJeNJnnmk3br0eZqw8XN/fbxEFmGUtolwQFdEcZS9k318gs0BrPNMp37ma2V3RlRXSCmXRK
Qp3qRafp7XZfqvbX2wuAQNAY6jAoiQPe6vAAN9fQPyjsiPNjpAu7tWRMZEwJMD92FEo6UOUjpG9v
dC1spZFxLAOHd8d52A+4GP1CpLNlOrDmPla2kdm4WH9Kfhl3OE5S1VnXu8bMEkpfj0DyuTJIoxY2
VIbBaR7AocLnk2Il83VYootDG3yWNmWPDGRcaeS3YhtN3RPojmDeDAYSqtdo99QwZ6smZznuROec
fDr6k1HuYokUh+STjKG2piwOOKUn+CWbz6AKyY+WRB5/CVzONm+pwnPA9nFUvuRYzwpI2ckC/thM
75h5ieCF7HoA4DQMHrENqhjzgFKdpxTb9Ua8XCXR9nPeg6XcRdy5iHlXiCJeIKpeIBsG/PKQv8Fk
tqzk3gkRAc8tzuovs2NMZ3/fgPap5LS6vmjbCdESU/nRoBrHWe5vg4exiMdRFxnt5o6ZAXCdPBCs
HBBNNd/wadXnkSQryMM7xa/IK2pLFFQrnNhmEWkApU7B+jxord0m930f1v+igdew0DztrL/Is1to
bDNFajZB7UhHCJhvuGTlgSu0rFP33npRNrGJfC9kC5usrBDXLp7kbg1ImWt4LyysS4mgFHD7V1H6
iUXtiQHBR9gMgu/VJtie8WEQqkLt0gJX8B8vB1F0ka2bYLbUjg6OKjo3eMHZIDKNQccvcJCS9Jez
XclgR2cPHEb8AkCh3BaKCEWxfCXtHypPGzh4Da+8AKwY39YvwLHfUvRgivpfE0iJL7UiYXYXwVQw
IBQO/ta3p2yvzXCrzpS0jP0378c4s9VO8t7U8pbXEJ0LO3vFV+cosG6j4ICQfB/10859NClow/aM
QuLMtgrmdu//iwnLo5Rom2mupSjTFOXve3PCf9YGPWCihBnIATm8l9VVRuXfwPDKb8N0w28DgZb9
p3oHOB1f/sgu727qNXVyyZ0MJ2W8ut9NJ5FfNDuiTwT8bW5SrJr7KmbkuSeGvoVYw40Ejnt4dWt+
sb3XkoBgPFkU/O8CmZmIDGKEB6Tjn+0AXVWk95p/ZwDqgnIL/+7FjB8wvapFnCaztrcuoMM+BW65
H/Pn/FqzNa1hrDo3M2nJoaC9k6Hp5D6Yt9PuxIbV2pXBeV/U++1qZMMf6sKGyrzxj6ra2LvvFWpG
JO+2P75nfNrRUnV+sch2BbvtVxhXzCiEuwDUOF63jfcxdxTzpTdc9QtAmnbVKOmvYJDQwgnBMGuc
T1c2c91hvVXB7UjXetJZdR0X1AT59BihZ4UXpn5HXp6ziY+mQJk7kDSUKS/L9I/0i+oUDv+FYgY+
ptImKyb41q2VZhh0eFfY5XLqeyjXNC9Ji0ocCcMDjfJwYdjqBmdrmBY2peloUEgG2tMpOT1d0PFq
+RY9IQ7NOQe885KtZuK/3KAVCfZG0qnfvmLRuqO2ATh6uVhCATXDaST6EqmZQX23Dixxqie92ksW
WaqGHuX0G1vIL4te95L+RIoSW7gQ28AFb1r+Ds2chOdarKsXjm7dg41w2RvjHmmAIammLMmQM4vm
yvvx1hjt8mzS8e+ncbNLfTSif/9AMzINwIhdpp42hx+GnuUooEpGK28RSCzb6CYK3PJazwBUFUTL
9wutQi9zGpOyKAydbi8jTgv9mfiu5rS1fPqcyGz/23W5dZETnBeFE1abWiMyKIQy4n8F7qXfzJU6
4yc3zh5fRG0wediWyo7o0Fm1YOX1AV7XhuDMWD8TLNnLsMJO1M3Gdk32X7sykPBWgOdc+A1uItre
p2OAQdQ9RTppKB9jWTRsZ4SHEjaN76WmEvG6RwmVGIInUhz8Pg+c5LtB57qtLjStW55Q59YoIDoW
tMhKbz2gTDPit+504PQysoZHx+dzyZcyNI4MDKB/5CET8HrfnkODZuQOPd9u38iB88cZpqVSOAoU
+30qCuC47dzL13K8ABJCu6YZDjXHtd9RKcyzA54wUCzn9VLOnzVFwAWlGlMtCpSQnqCLztDPM3b2
K8cSvtBN5f2sRhDwt9oknah08/ZiyuIyp0r7XsVd1ma0bDpBMLJ+l/4Mkd279liSJStgHmVdXiPD
bFaeFIwcQu8b5auF9x1avt2BkF5hXas5A0ZP0IW52JMlUDGrXZBmlbpGXmwsv8b0KfD995rjugty
RlEtaC+N8fpPSbvJoo4EN8StjAiRuqqqATk9FaIITp9W8fEacN5yVViQc1XI7PlPPARRk9Fk38zA
TO3ZmJjrqjDALK5rwYfQmhm4JgPFdBC1LnrMDJW3M/K3JR2oSRAzXKI5t/8IVtNtgVJAlM9V/6X9
uVpfj75znPsqyawNaGIJuGtngvVHqc4ALi1gxEDB0gDiVz6U1F4SPPKxbAl5GUccTeLBHhZj91lr
R3DqxuqYNgGVu2SMr7Jr8domofleK3+N9DGQ6BacjkD77MAlERuwq2TN+KLyhBEsMes2zbI14XYJ
GHjMDR0hH/ScpAYn7sY3h3ylrJ4ggRbvuhnOZvd0BTrfEeWhWxrRuOG8Qb4CrUWObZWlkKanK3BG
jKJHim+bqaWG4W5Ya1xA9RileT6Wkbw/V7DtF8K8ZD8WNiDh31/e53DreVgEy6A1zu6XWtPKk+ow
ykLfmA7lRD5HAut4/3HsOGlUurlXnno+J0btH30EpT5olGmUvns0Gmnu3YeJg6TO5/Q5Sb/DmkzB
xMBl+jk9rBHI26cMmL71wrL2K4l7eetr267owWFXmmizmgdowE5vrzDhQzfMAQvb2z9tNfim/HtJ
PITab/k+J8rUYbW54CttNnFKMZkoFZfVkLdqD9NEKUl4LK9OVfJ7RNlY3sUWXZoCXlEZE7RtTueE
SRm+HY+UsyNWNsCP/QvGAUt77u7mAXeqpml+/oviyw79p61DrGo/NbVz2uBHq3mterGqpMhskUqN
cE9SnXV0hoGgsrdnmWl5PP3Gj1fi12fiZbeEAKLZGQVeETLvh3MsPZ3X/KzeR5fDWJ1S5ais8XR9
2oLBVjGGfizNc5FUdNvtNonjetj/FZ7/t7QNoqf/Qx7o38HXwBxKR+LUxYYr3L17aPT2f2qZ7E2R
AQ3CD/U4dY0SxjEbYGnnoZY9J0GxqwR529Hy1uXOopdO0nUo9zr8QIaklyg/hjo46/84eA6w44YQ
Qt9JW94CUSAUGZ1eSjSa4HAEfGraPTtK9ZbEZhfnlkDNBz8+1CxTAP/coUuk7fZCdtJIRVKxn3AR
p+LW9lwAy+GNfGwliKAM64YkhxLMGof43UPp0EEcI+8/5ov4rHQBiZWbglRStT468kGFn9ojzoCJ
t3ApltoXKUZwNRhLYG55DQ+fvdwZM0iDhGzlEOsm9jDPTGS0GoXYCh29PK1D/8TuphTPuPR1N3Pj
LoGTxenAY93LWgCBwxPBHRRMuJtcg+SU0VIrh2stxI669R5nmTnmuNTQimytD8ZpeGVX2+Ffh16Q
HZXl3hPaeynwQ16VheRfIdxpPftHIFV+EKwGE8fz7U0cORZQkSl3K/lBBN/MqNdKltOETOu4fr1F
Vf3ovkFYd9GYFO6VD4G2Q46KQV/eKlZvcBH8BtzIsjs3reLjthPuokKXa1CDk7XzLZXwe0en8g/b
4psCbFRA+Bo5r/z8jZCoN0g/nCk+DjrmQqry0QiQTh+uMISLHhDj263IUuGPaUc69byFL3XS8/o9
sQ4zYIkQkoFTwfTY5QmaSJqHjSjRoAr2Mvw4Pa8IGYAZLkSY87wLdnKYlsy3xRrkKX/oMtgw0Xes
3+FzVG4seFIvljXNqwPxJWxZ8I+loavQaYBPTtdtYclSCVCvk21g07JJzBcYaoa5k2HBsQOEOxG9
EsWzKCVi92KlBQ/f4r1oDn7clW1V3l54t7qyluPBqRTwGPHFtGg0ehWmCKOb2NdQt53VNeZZpLuH
qnEWvEhHpSSxDjvt6ftOMq356fNxfxrR1d9qpW24DFV/9s3c2fqfh88pnb3nMS1T9eiFqGv//4gK
rZJqwMfk5IL37cmVQom04WKgjR0IgQrGJ2ScArHD3tLLpkSMq0IRiyeckdaylaHMzgO6AvZFZyVS
1X8G3ISX8PtGdxjeVbeoopGU+RhPPpTDS+PwoDBf7VxRBPupGw9CgKVXowkUzoGxA3SXpzyg3ya7
ZhWTbBVU6x8TxQimg77t2F5uHIW7A5hh4/aMMb6tGYMGOmB4TjKCc9h+jcgTt+LaOM0QEXqzHO77
NImG0/P8mUE3UK97oGcoGNByaxEUYbGMh0h1CD6xgjuQQfUBCI9J+mUt0iyOZjMYo4YkqYI4wiw2
xEO2Y+H+QGlGEVoBfQtlKsyX3Lp0575wu4TWye5FYDMIafOWOPxl39rof+zXTvtaNITJyzZUlTEw
mAXrZ2oDkuR/DnXyF7+0VXJmpV2Nz3ckNwpOd9UwLdCLa5smzlEQAGZpqf7KwDQEHE0C7oA6uAbC
fjq/6UVqWpKVugOOnIlk8KEAT63FUlhUOiTrka4aWcx+UUsm1ykWvFi6FL8th8YkKyPeabsrQXbR
9VrWQr5eJJtiudTevmw903ClOppEs55+9E/3PPEqFJ2AJuXk1jz8AoY7KYhqR/m7hFePhzNx9+Ft
xvorAvz5JGOByyz8c1ltk+uxgrFv3sb7JyQrSeWOoEV8//vcVpbmWy2EWPDz1//MsdvM4O7zGclA
3tpSCGaVWzrb4hpGPMOTqcyBSO7cL1l9ehx1u1AjF9ILY9wmUc6Af8qKP9fylw4lb643UVxfq6/T
KPBWrl5Ec+YhVqK5yxg0+XQOozRbmiD2Dvu5LlP9hiJImeH58qM6xrCf8D9TgcvbhZL5Hijg1PX4
sqFK5Yed7ZEjjTvvGUzbktiyn55NVpSrHbUnPgNJCHn1cSPWAYFjYXMiz2598FhQsB3zamEbbHSH
SnkNCGY2bK5lmVFmNZV2EpYytL1F3Q/HXb4IgoD6S66zFgareNF4nRLtPP+JfHgQZ0covf33HQNe
uLoGNQEZXXnEXLrhKiDJDKmuCh/dA4AP0yHNAjpBHH4xuzCS3uvMQliMPLCohnVSadtMqTY1B5lx
S2WQM4TdkXUvJYE9/ycOI5eXGutgRgXXYOv8t3lj4V89rAaDgRv7oLkySy91OIAYQOvnaau8xaIx
2UYsZs2NZG6Kg03+5y8SjIqkgWcCwgWFpsDn0WrztKDnLZPH9U5SQOSbDJnvILxQna8ZJrq7v64P
AE9EUKkzEhEF17UwYW3DqBwB6CibdE7mLTozylQPo9F41i8itMmE7jKBi4ENdPJN5AU4c/ADHrsG
jmem1q0t/RVqoHmOf8inrCxa5PUXOKjDgvvay76EZPMgr8BunJ3eBgfB9OjxKJNZdHGBEkL2ZzDo
lkR2ofseYHSQKtFbDX51DdnjUOT+CtVC8hdepMHeTusKd4AbWkbF42WYejg/Y8WFLfVdebqhE9yI
f3gHJQ1ZdTuHmwb7Zqk2QClala8LaIOcNg0lH3UvHdpN+zMQ8FHWAFejmHdeA0iWpol8CKvWeivs
3ykKl3WyexdhzM0TkMKyrYqJiSkBgn/zYmpBjeI5iiMLwnf1qT3MMJyvlGzbEItzsHudm0KH19R5
wyaglLSSKBR5+Cbqd3EjlSqysyQgyABBBat+BVKgk/3p+Qz3y1QVsXkWVeZLKfgShQIzBWQlRwmV
fkuJ2hwCA5IJPr6PVsorBCsKx3VUHzcIyr0f0Qj/pIGzm9ZjvuhQyrVCrAuc00uW/V0BngVfUa7U
eHCMDAA3vAQxj03NmJD7S79uGUBhjT/t6CqlU5MvYn5kK1Y9dqxIbrgKRNK8UjYGqIsiKM35lY2e
FucZvVPI6j/dnCPxWo/UESrTR3if7F92XykUFH4ZuG+Gp1nUjMxMsi7eN7usFHpJ+zfjfvCnsAhW
vsmsYwgCRFsFdnnFRr1+RWYiiKR3QtUG23Bjpe2tATKptaTVbPVn+pw+FuMg7ercnzh+QoGe+dK3
iBamg0+GZBAnZ71GuDvYQPMCwi78Kg0JN6QdaeEQ1jnHGOjcCIVEhc1lPjpI8kEhNFcMMMbXXfXI
TqE/iQ9gdQwu+msIgSgoFmMKMo8fTxdQJPMQ8928WTXZmNqQDLmUnLxwS7y0OnDeSASKgYaa42C8
L7qI4zWvK5wqlEYYjJJ8qS/QaybIvO4PXpdb+Ec7oJvnfcmdGAhWM8cFP2MfvuUaA6KDYGwD3rft
NJziYF4sZPtsP6XNLI1PDZFWOoxX+sEIYV0mMzJwbzx6FP0M2m0bRmMz08cg+PvIO2IMkQP+ejGq
09fFDF/XdRR2WoXBGhoocSs5a6qTHTwApN0b6RP+zir1hMeqSPoiWUWE/rMl09badtRJ6PV+EkEU
cQz/1ZgrasBc+CT0ptCHgJ4TNLEJwD1ci8fwm5HmPWc33+A3XN/NYG2sZ4GVDzCVBi+wML7COkgx
hyk7yN37UHpj4h93tBajCqU2HsJLF3ntgvcbzSV0IUx/TGo29ih3kPxEOajKHBdffGHJOwcILUy9
qbXHbthuoItWLJQCfw+XO5VxxuyDbNlir9SZg35oQAOd9OJMKdGMdKaWAFALBAjysAcnbTXWtq2s
5UaJWVCcUhvdWdrBjgQOWvjIHD4xMDNUm0vSvohS49fGKWp8EDjFE2NJt17MBebstuhnM6KhMasf
YBECboIrBF+ioea+RTIB6J9e8hlGhQCI5l83lj3GyGb7a0jsXPRDf2MzDlibR5QGngODy9Sc6z0M
0QqY7nNBFIrGACH5cy30bivdtjgjhPYys8fiaQv/0rOg9jWYsODOl+vltCW/iJsAOR9rm+jGVrf/
tonlvzgr33R1u2TIOJGvVjUEb8zk2W1celBdB8H2J0KnFxlP8+Qzm7XUeQZz0qtBN3h135+qssGY
MzUX1ObXVChu8pGvYGzmuPEu1Br7V8/9G/d7UrFK/CDF6/hoZBwxH8wWTBLrJorzkiinqg+Oh1Wa
QVZY5q9dDk4JYAMy+H/WhJNA4sruShKYiu8ieWavLDAQWo/GFTrfIowCNY/GTJfRiOZzErpMGkYG
QC+JrbircmZ2fL0JmlRXi4osW6w42q2XUbN520a5CbO9umITXiGqPSNL9GuLUjTHhHlHnqYOYagM
Q/NhVFOsb0lb2208aHUrj7tmpfpaWrOYZumSiZ04OzCabUEM5aQXwLFT6385uAy8O2Ygn3YMOZco
dwbaf4+OhZ22pp11QZmuTcUZ5CKiuDEd+KvyFqwrampFOLxCMPEIJ8FfLgJWDgytsbhfi/4rvIDi
QM1LM2KaHJpF78Y/JYaFsygO129rrmmMu0nUebSQvCqt1gC5PsiVQ5SstcXeggD0TKWedraCznQw
vgtkl8iL6hJ+mVoXPFqWV1ykVVoHrQ4LSXvg1zog/kvkgz+e/mHPynR70M1c9OREWpZJ54Zpw0D3
Yn/UdtkgRS3Eo+/4j3KaMapzVOpAPEKjvQ7IaN4KEil/E2nbBKxGkMR7eHDBPglJFA8dSzo/WRrq
ugB9+H5vtL3R9+Z5tbc7RcvCEao8wjUsRPxNeWeBtS8NOtNfCK1tFFIwCH9JZ4piIXJzZtQBdabw
0p4KSRVf4GCKtliOQLOuIAtNmqgdFShfrDDmp0KnwtY/TZiH5q3DlhPhDdji/igsWxP3PqaYY07s
voLTZTK08qh5pxSaEnH8JHJ2b/WOP7agfFH/HMtU6aE/qpHBzMUslXN5178GknyQlVKBuqQQcT4c
N+CHYqdyXUgKH9WX9heips7ljR/rNrMwVgses2p+QdNQQFT30z4STHdXdZ7+olZw9f5NHdoJLvbl
OoBWndDoJApPnSXOFTynRN7r2c3oiOkP9Kf6olLagL3c4cby6/LtXmjm7vw9wzxfDhjaLiRHlAWK
tZ13PNTGCCO+Ji80fl2T+i1v/9ynoclwGhCel1CAXs0eqG7njx7LF9AWKEqgkWOn/3hLWcvJnm6d
554rM6A7JYZoXkreNdXN7nEguRYEeSS6QsFUgeUKKLSiPZ65bT1eJSlI2rakTpjZ1eluW2jX9lb5
/dt40g6oZX2yi+wZsuTrvQ2Q1M/WxiwfJz4rU88YReM3erthAkmGGFrxxzYzCzCIS81HOMZgdjzG
6p33fcs3k37TtkLr7Sex7mdhoyZpbqYyL5Pm+aNjOIL5Jl7BCKIh6QxhGe0Yp/S/ZhaB8nBCzQco
5MAihSI/VsRiAVY4eshVGRNaPEAh5xqkd5yLP6cNYfL1g6evBdyPZ0dgGK3BXi9JVbkx4nL/ol7X
yx/r/7fHhwyKJUg0SPXPnTc0bqqFUgia70Birgzlmlq9HS/lUQDxNOpMSBki40nykUelaN9Rtp1d
K76a+Yp0W0WYmkfI+Gs3uTn0DGCe6umu5VYcgnnRBky/SHCFI6Ft5rrsNqtfHdzHFHJvjO7lcWX/
FfcDtDT2TWjoHwfCf8+6RmMzaki8t05H4ZPguD5PjqRPYG5gxePKMF5E41PZ+VTWSC6HTsqZe2J1
oXaeyeCbh7Pnkf1BKPcfNh7UwWMHNlCrk33hlrhEVNTTxF86SkovT/9youb4+Fi8BOrjAjJwJoTX
U8utMJaLg/sC4GX4As0QaI9fDPdFNCHes6mZx2MD1aIIaL6nlo78En7YxjJNrUWWnFrURZ4cTHFO
hFcslaKnCnV1hiJ7LT+NQTijQNdUI7DM+dW31vo7v7J3VKwoBHTGJb22/qFXHcc2AJmlESSUL4gK
1B2WTfBq4kCTee89u3cq7CItyhg38SVvy82b7BlBuIC+psdtmE821g9fUoqEM3bukcS5vMFaT1U8
KiQXfKmmhztliou5kCVGBqm651mA2ynI/BFyrClI2tooPKifKvJCrRHNavrAlTxnLm2frIW7/gtR
ElcOGy0XPDQ0AWMXlBvRj+wD0tfBWtwQted/GLUzssBhVQess0JIkO513m06YynkInVt79xjOWAc
ysu/s94vERMCsrOEzHkSPYHyWA8hlwpCJfaSJsE1K6L7bEc8uyzePV3KwD7w/RpDkdFYH3zopXu2
xVQsCSjW4CCM3ss9YCHQM3hgWxLWXLDz6fnl/iYo8mUf/fHbPl56j/fZ2xc+AijfhQ5Sp46m2Gwg
o/dlYgqJVeLFdRxDUIgGDcbLT4XMqCHcJeIFDUlX/KldVDnM/wTOJViBUDxJFI3KkTiQeGTW8fi3
2i1jWPnEptdYBIqKx5irorQhXs4kL7xHkPs5vSg9Jx5ap8GZgtwZ03dew2f74E4yPTHIqzMjlvOJ
Uvncf9GXSq1rjURcyV1TKkgvHYUjV4AGqzh/+cL/J1H2ECywQLmsvmqxUEIw1nJM9/eL3mtV93u8
5BiuOlzp3eAfmKwH5At9Im9VLORCPbY4krVVzfZZI2UHT7TkiIrPiT+Ph4x/VQgx3w1m5cWJblCm
E38O+Gqi4RRO2mIlYmbLXCEF0cdOuc3BNJoZoHyMWCSAU7Vv2kt8IPgPxPXcnW44hysFXNfZKG1t
KY5AL6uaxwEiExbxg7/j6vVd3hMVrM+N86OpYtjpp3pPtEYzl+XP1VLmmtUAYL+atxGa5ixXiQ6R
Kg4vbqORvMVUaRplh9t/WRhI3rhcOF8OrEcDW11EfUrMIcbojMe0k1TuR7MMLiDEfzOFsby6sVXb
NNU0mESez68KBOa6/eWSx9qeEp9EFxZLzpjRg4aFJO5LOPHdlXqk7eDl+TvyvvRroRI0nJ40MjTH
mn6up/xYsugaRfWxraBuT551T+VlplTwFs4gecogH0x0jyNA9fLa/xQjkSlxvUBp4AMuBZGo8jLK
C/MaegndLX2URzoddzaDBzbB4lHS8evkUjKhw5ZZGKmxPVuM6dA9W89ck/9YITtAFg62eCnu31Su
cCwOFOC+q+LhUCuXzLiEE88Y/XrzuMa12URYMtL0+GYLQ5FA7Gi4+5MGmyBfUlnnPoMKoyj8yAxu
xcljQjnib338z9t4g567VQCevrPWJLRitPM8dNrGrvk8y+EMpQ0raWj1i6AkwcJF+OFJ3IW/OS3/
giDrbZMpX6aVhcwBxIqgH68Mk/hvtLKsRjV2pFmDR8jiOjk+wcTJMhWpWzjOet8w/SNTWnPGYft3
xTuCHtHTxaAJRyHl3D9o1T75UyPgr7xVbwHvEGgAJxJJRjlFewX6fllyQTbCoqOGsAtAz6fQwUEg
P9XH2GN2WnJenWNabNCzjh7k6MI88/4bVCxpPBJTyMesD25bqeDUkDHOB1q072zHHbdFWlXhwH2a
ad6Ziv3Im6TZOFxeN7G7+7mYztb5YkJUeq1x+GqIdvKMn6SyLHnRIRXfUK/wTmzyqGpIw3AF5R3O
x495CASV/3waYkgkUmwAKot1xFyt9lotlDsSNt8J5NISvLQ6d2sN8xfyNWJGF9eTnWN5T7lSOxwA
PHZ+AlLfvlKxotzKkZXcTWNdtCtoBAwOP7o9vzPdMRf77o+Yy41b4EvA61LXJnPtWPOdDPS7sdOM
VnFAEtcHbKqk5BMXqPgtoMiZHakatBaikI3bA30HeX5eJSHICllCveYkkW+CkBy9ockt9kq3wUOk
tTcnG9NG4nMbaCtmE3Ws+hbDEt5Kie5l5rFkmvWCxU/Busw6mgyfl4WkPgOmOnx8pwxrnrmCQrvV
tWzVuVPu2aAeXLSl8+JvglXYk9KqprqTFqMM2/w93oKeH1cBSW8pFv4YRzBnOiaKgoqOb+xPnRHV
CwRY2KSO8fCeeQ0TYBrEAUeIAuRM7fzGP+EAGKKmBO6S+1VuKzgLxyC/YzosaKm4E9WVYoKSl8dL
8d0+fpxYp+BAoMRsVlhKGFCvXLBIrFtE1BWZkdT5c+SLQCx6ir4eP8g0ZnR44Tn4mHggNbmclHW1
3OGD+30mvDKkJc2YzXv1hqe68DFmS6IDzRxsCQXu+dXKsVy3CXP8IqH2Vv+l9T6h3MAQfw7fHk0P
rUWrKrbQQf4qOH9BitV1Yj/s2t2+/6S/qwJptKnYwKBbPZhjYXktr+mcr7ommBJcSsvJLfq1OVy5
/ppwIgLMeI0cIrGwdS2ajJnRpiGFOXhgYoodMxnIVa+6AlYJKfhyCOFYUXEshJsQjLf1pDTz7OKf
YnYXmCU/KCgsJ+SBuysc1/EGKmZz7WzOWG68rglWbv1rJVu5TBxVDq7BPjl0nrs3hyCWvlmN8cfe
GfC7LGVe6FgXLrufczyBFHXlgNRpbHm8EHpgKFPU+I5cr3PtM8H0pOr4JWqbUjNxhEuECcmMlf93
r9e/q9lB6J0uxziQH5Zf6LFwOsfJfnP+6i6t31f0uBJeAKj/4NhzZMi2FyDUMP8ED1hTw2EPt9Ff
436Gphd7Lo2yy2bmseS+fSuRtqPSJjj9SLaQpc0HY3PXxTfzpjX09aKpaVT1to5SSXWUs63iwHEN
Mf5v+PLVQdHsqKlevldLWItYA63WaLcbsoFGfdHdzO1qpUkhHlSdG9lBX2kKh3QbXTK6C/WiZArm
up6NDGxftI7hK/4u+Tq+MtenrXtpiIrR4lGvN5QcQRLIFtuX5oFcOCtQUZQkhbocsINFfGxU1u5K
miSAtBhQn14LiHNyHci91gnBJHoFRpjhoLHZiqU3wVDrZScme/1rdOl3AQTIEwy9k/W4zZpEzU0D
pfa2g6NssnvxQcBL2o5EyfRsaHj/T3T3uHXtNUG0klM+9JJCrgb8c0930PtUh7ukjOLIeKqhSvD6
qcll9e3LbdyMFI2LPIu0yYLdTyZqqjstniy8b345oHX1a38COlue66KeOQRUF/ryFvcssfMZFejv
JNXesPU/Hm8dxQQAjaHbcWQfZ1oRuJ3GaW3jxL/3OS2z8iaFO01Gq5m7uLjzXJBFiYMJ5lRkG2Kk
WN9kSzYgDU2HRE+HGv1JXcrBoUMmBZYaY/XGHX4jClSmueIZu6/DSut9sRjw8565rD6il+cyso/R
gLYkgnuPUxKYoIlqltVUYxUlqlETQwU9dDyBfN08P52DDR3sAeZ3Ok9NY+Ga/hR+6r3yNdwwWUVO
FMdI0zEpPS9UwU/p9qyB3iBj+xbNkvzYLV/Z9OuSkn9XD/tJ2iYB7h1Fx656qBtwGz3gj06TEKgj
Kz8/qHKTmjrnV8OAWjfGqmnUDCc3KVzI4r682XXooheEXpENK8WVK4cwFksC8NwP9AeUrIEjqecA
Fpi9GnAcVjl04d3lo3GYxs9ZPh6839VZ95p+TmzjXi3wgScKcNyGAeGIozYjCy1rpXX/abfWAS57
VRqM7FKkkvAHd4+0rZu1YURve47OEkghTKkL0G5M7CrTz4uYQ0KMYR5gInMrq16dtpXG5VsyB7K+
eiciXKDjK0edkO/I+gCre2KTpk8yzzxR7EYv2Fx9vIfXUogU6Xjn5jSHNvyv4tP4VJmaXTaAS3JM
+wBBNJcWK7goew7xaxSFrkA97Yb6rjtNDGooHAcTKFWf+iewbKEpxanJUw2vkEkrqgDZvwgAQn2c
Q70+YnNPWvk0aWo4jXEPn6xUtnQYRIWNQHHG+UoTkzbsw4ocE4sDG9ezTN3duOqprYz8cxE1jGAZ
iS2wYBALKk3N/z/N0ba7ghjhG3G5rDrgbLEJDqY7UPMTrh6qEmdMwnTzl0n86QAvyhC91yQySzPG
OmH9XdK/Azp5IrYlPBPgPqzJ6sNhpnWZJnMCahxLTraDviU5OZ0urCQwvcGUyaNnrFSkN97QoSh2
lgz2/JWFxOgWqCyP40Pz26yyRAVw/orzbWgGKvT/v+aY3JgcvZ5bOkVbgiW3ahQISk80jSzG8ELh
8gfVNRKndydUJQ+QtDNhqtcUpwLURwmoH1f4NRgbtWY+MgTxdCN6dVTKTQuVhOASrwQ3S5kS/5Bf
o+GCE8vcFmxJVhxdvTyEHzusAfUh5AcjFGW3K/jzPsJYmE/CX7G/PkYzUFCTc08uO+cKDUsj3/rO
m32noxu/QEJZVCAyJ6Ev+gb9tygULYwOCWQn3pn1blOWncZsptAI+xxKIQX9fUXJV+FzqC2F4ceH
+HssStHj7cOTDOkvv93Wc5ZMiclKkB2PQg15G2KE+DNf0C2IaO0aXnUnAXZrlH5MFtOCQKhgbPei
wD6VVE7BCK8EYv+eXAyZB3DTUr1ct+WDzoHHbt1HVXKRKXVeLPRj4+wxGEh9rAiDY0bdJ901/dzQ
2KiQweNQwy6furH68G9hQTmO44yxaDz7XytI137xSlT6XS4YotsGphSOkHaGVno68M5iIjSNvmia
k52c6xbLblqcRJFvsJo5OMEOn2RgNroE7KBQQsDmcNsO4poWtwX36WPRcm3RLY64AXgpDkYb+DHL
H+88+pqntn0BGbemTiGE3VsSu9aFmZFibju9rNZsmbcrvRqgL444K+e91tBbwADeDnQ5KVShUhTl
IMXQwxqUIkppB1oGv0l/p3G7yBZ7H++Wa9dBjDK4P6jMjKtDjvOIOzUAtMO3gL1FhjBGI9lFgrTW
uoouAKpADlbUybPeXMtoX95jfsjmvlqRtpTxuwb7Hd30uw9IZi7z2vChSlgHGuKdgNzo/XS0MpEX
6NdKq4qEAiCdn7bmTf+NRtGyuYRH5lyiy1+ojPQKvNJgAaTno0lqB1S09DYpzMpklaf7H3mHAf7c
dEU8tFe0bn1v3RfxRfqKBPMcdV0LqFvOzz4lbgIhkUVrJIXxohMZk9eQaN/FgFh5mrwl4TwLUdWY
RRnHJTMjJzo3Oo+83J3DE/pK8xFy0u4dFLapHJ+Y/vaK4Ym/TI3+pco2/8E4B+AYZrqcAk8bs/tt
OHp8TNrd+Kd5nYvKpU73g7lmNhqnMb3j7yz+uwNWbBPIqDzkivIoD26vVQ+O6hcD7tHt5SOuGT2i
Js8psj0+z4aFs7wpvXSCkikah8c14BYoq3GT40XHiczyZv7yjYRB8qVW2X4GfQG0NIQzky2xYiS9
duR4hSshv7r3j8se0q/Pc7eNvsp34oPhltlhAntUHkS0hhgpDjxfBl0tdX8zi7OEsKC/sOBltYdw
QkTg3sUJ6sL+1oW5kZccVCJR/8LB0pFfT2AhTk3ZXTBrt7n9yPtntT8Lx6zygLgjrrCj6vmyoocu
R6GBTo3CVm/CxLcTYh4bHcCVA2nvQqzuOV/fENs6XgH33WmswG3Cce5jMHNNVKyg+bxuJAkGRKJc
1R0q3bRkoLph2DXGwr34NdmCqqjzUwl61KqXitgZ32g9dKp8ngZ80jq52hOQVj9X3lHhfztI5eiU
aIOqohqNiOVbVz5GDWQyOG3l16bBA5d/tHhGBcP97AITP00PbYUOpa0UrQMXFDtY50Rxd1lSULc8
KAoIPL1vIcvDueAeiOUbk7fZ6/C3+LsIRjYaiOWycxWzBUGnATTF3ObHi9gDI1aPV7EUb+p5GsLz
9TW4onwDH+gldTn+gFYkBXdS1/tW69kekvSE9tVW3dtPQIpTg9bj5/JtP+l//5VxnArIo6yyjhs/
aCbkF4S3TXGhxSNnJ0iUa/G6y4pncy8ViJq4eCy3yHskcDnSSMfe4vCh43CUSaQNlECFKalA2XkS
ea5/yhwSn3obRQxlqZdQ4oNmH8WhpF5Vo+gjUWAgQdEuPBJicDKbvlPftkE7dqNn4kMo9wXIslpI
ARjcC02kRfyrpvEyZdxHD/mZzHe8irA0x1yiTzaDDk2B8RSqCl8nJVpgMAVJxFcduICmCpK/CFu9
TWhbyyJLdifx08yN/TfwYMl0OaP9oevF/FyppqvDKCasGd2vDhG6Dw5C+jDL7GNIwOAm08N1YxSw
CAd3nzmycyLs9IbnjjGcE3ssEazm2GJ20HTPArQDTN0LlEHpPSBZcnSnVeOlNr3wfkAOSDYALMuq
XE1qvkR00Swi3bmMR0fx+burfDA4W74veh+pKXWo3X6TRcJCOA6cpFFWVcCzgIpdgQa8RyrgcDG2
wUAoDwIzBkdRlWjpxw3I1A0Iqx12ApjS126+e7NXhkgzoX5yORun2YnoWbTnLtWCfxDYKUn4kexV
ZSVvLj1mWNhzc4frxfZpcxZY9XAgvjJ2H/Ku0XN79FYKNycnWdOu780uyU/9zt58I2V2+QgPOTto
dVtyLKgnPQLmYuMv6hmUIGrK+FvEFdPzwhMqhcrNqezdzL+LWUA2z8mbYun6w5R6DA96Y1f+NIwR
L4aOqfA3NjcvCZPK8oE4HYg3EJ1fhfVkmsA9MWhbxstg0YEtNcPc6Ujkh58gPAL+yhSaTJhEu90h
dc1SBZnfNfp4TW52W1OUliQQHl8kdhj4yMyZRFGEpxWCT/HR/iirR8cgI76B5kyAoj2t0qhn4G9a
Dk76QcWYDKuuRRYH4y/CE8Sn50ibx9euKp3L2V5xHLGI/mUtAOBcn4mKmZbSbAG1qU8z/hd8Qq0D
6m9IK/HXMefdNm/anT/YOmfxhRqbjsoAytm+c15TfMYzVZf0ZCgTGsQ4IApY201DeFkvDm4ldWn7
xHC006a/Yq6JkJ82Dd1XN65K2384eOt02VfEAgJ1y4KPkGsEGbZemqFKVa/OIVnxYi4ZsUprulUK
iNogsOzeuc5cNUhfQ2qbNhOaVC4cmGVMuVnV3d6sQLcKQ3rSjLzk2Ndly/20NyDrXoawMC6QGJRh
TAkolANsjDQG0kC6+rITSxOdoRr/9I4FUBZk7sxO4RVl7iRh90wijkPz7qgsREqtFYyXXzRiJ7Vw
C8eHA/zs8jZg0ImJKm/91M8aMJO5wsm7WhPrMMAs11tK8Oq/g8gB0I2pafXaT01pXkUdRWHhDUDA
+enCWfFjOKVujSWP8Ou8AbyLTKoDFuxKQDt7+gkcceHoT2gnhlo0YD4SU29cVJ2CnB+DPNOn14Gp
ix8beh+J4pDdzv0Gpsg3XazMkl20q58/kWgw55UAXUZWKqAEw99uviqClzd7+OvceNmHFU2mKdZF
sxwFiSRk7oZncKAwATWI6QSG11yduah4qled3J1h7gtMnKJX4LKwMF06dE9oDKlznAuYOSmrIBpM
K+ORv/fbKaRIvt4pKDZOaTsQFsGVgnxFc5MzKmre+uR6xz7Rx5EdeJssPUtith7zQDxQWGhL/Fzb
GwSxirOP7GkAYi0OYJXYPejZUx5B9V3XPtTsWjVQUErOwrXdDt1sHU3fzmyvVLT/Kbpi7yll82PN
Fsv/dNEKXuwuGpviNJ67onIsfEkQoANcyCo7ArLuoQGLZ5hs4SYkxFz9VfTGRBuD820vK2oASZAB
Z6wi7JrRzCdlxlNijKRs/wjpBwk849nJhIYbdJK7e95AWYDGTVkcBSnj6MzqInKij+CJR/aLidlo
ki92Na77PKJNrDU7tb3g6lKsb8Kq3SGNFeB7xIUu4o2jqFYD7PnUMh7Mdqh5bysj0sH42vmJjc4G
tAzqcRMrqf/B3f6KBzTJ7k+YeRF+Go8oDwudp2eEDbIxRgI90GnMJksoxpoumo/U7IcAhBGMK3xp
lzBuzlcJebT7+UjmuyYoif23HhneaL/hdgD/HqePScC4mb2XR7mMdl97kEPVF7Fg+OwX135UbVMg
CXhittL7X3rHXd/sVIu41TnyRMlnDwJ/S6idfpNTnZ8izIqaNr0OF8r7qENvYTja/QUKuRuJTkbY
koAKt8yt9AwtzKDB/xqbgVIqXqoQwkVVu+27uSL/POW3pB1Esm9aBVZz9P45mzf75lZvQzAop4Is
FQeHsH1ItrK5WTKdeySCGFfVs7yF0qEIzqDqxMdtCgyjuBNCM/v+1bDJqfniDci8T9XSIiBFGEkE
JJqJrRU89V4HpcGSn2J7GQ4LwA49eaXJwuigzy6Gykcly2QXWV3tw4LCsOXESuTHRmEIHDDwnoo8
ZvfzNH5Zhjx3zjdddQp+CP8a/qriGD5ctsrneBwnwyrg6P3kLAftj+Wf4+N4mqoGEIwknWKD9nTj
3em3399J58s2qJLX1KwLlUlvqbvuv9iWAQh4zl5Ep2F4Gncm9ACu7Tev5yIvGtaXN6BUcqVI0szx
1U0Mw1aHqJcph4ndpO0YEsxPnN+21Pcblc6nhfwzW7a4YGlhj1JqGPWBBYlY0fuUwJnmmnH/jrLy
6NOlHtcd4FzLPpGFbvc+QU0ubMwCOEkJYjjpIKxlouzDoE2iWfmjZ2XSfjN2wN7wM/12RTHlr8qW
3eD8upfc/gAAqKvH9FTGY++1OI89cWzfo+0KHA2OAUqzCswB6OsooDwHh6WjgWGT/MthTNqrRAkc
Ky+wukOHATJg1NIwvDwp8cn1YAG5v/AcBnLU5tIf0E9FlbZ1e/F7OwIicxjiOzPZ8PVBx9KA5pAb
7u3VY3bhV0VLBBza4PEATVjEx8tInSLcsy+0FFq9vHpqS5c7paQA0TkBGYJnYvDja5/nHpx2WqPX
QOzy3zeTM2UoO/Nq/Cn5RGjWgS8b5t8aT5Qn8oBP8V67xRCTNnftPGahxOmAgO075jy0j9kAP5Tu
/fwNWEzsZxXXucCd7Di7/HAsat/YtxdqMjU/G3gGX0358+Fv0ou2+wLIVkDE/2i9n5aKBX3F+ccL
7YIYb0YQLwt7LkLw+ehNmGbNQbc7uluNp0KN0GtUrSlRXZb60h/oFe6c2ewU4icS2MaYHZxIpGTL
dfFKkyrFYa4c5bvY4k642IEECZ4dLAztTfa/Agde3Lb3M42kA9IehYiVfvq5wF++43VYBSQjahHg
hdXBGTLn+TcfBDV5uRs4iOPGWjvK+lARAB6/EQ3L/gsB9H+NCLyy60nXvf3/u8gwQy6VHASa1yNy
ikEcxmUooRP4YgXqSC5fUMoLEJm7WNgSxDk2Y5m18Sg6vaP590oBSQ5Tx388LpM/4nCgk93lN47o
NIZfSSMcTv49wWUYJ/b1Du9fLBn/CUjTfNgB/DRABeEQucHJ1i9wm22KIk+IYJMFKVVXW5mnARjQ
RucnZIBP9kONyqwGql5yKCye3TMbf5O3Ddwt2REyb4AEA1qLg1V5PLNgare+DGXQCabPuXNaube0
1jqIlubADrCj1HIKFUf7Z04xv1Fd8kkhqJQRfieSCQhOFMSYDYYS+GrvysuH6QukdEsJBmzYx2IZ
HVQp9n2tURSZfU7ISrSZk/jO8nh61e/ykGSMMPsozL30Y1oqLqr7/4n7p2i7pzKTpibPUIKTTbFv
6GrIsFmMxDvRPQat6nNpE6yaSEt/4lJQ6LyCDK/MG0gj362iiOVMhzpZ7l+5xN9SPBGWzFgbP1SJ
EGSa2gY0jHLdVDzVlKBwIS2njKRduASRmMhTSXQ6rrOikIGvy2u5CyoKhEgkaqs9XrEJPwDu6Ufv
JoAlYPNDFABotP7R3m+BGxMb5qqN0u1BYBVkMHWlfdV9s8DJNzbq2wpiKU0q0P310zBOPfdKDEXm
fqfwmVs8pTRqu1VsmAY6u/gGOSJZevod8Co11dgICGWfrpZcbroMuYvO0eKJMwbDnb0SesoibcRd
xpY7WUZ/EnBD3+xqpj5uMzPEJ71euAU8HXioIoKAfhHWoR0exDjAntNa92bSPXCtYAkEkZ8KHern
qSidxkhVuSQuJu+UcgeG9jGlZjEeM3ER/EcL2m60IV4eSvcttx+4ucDM4fWrBTCQnM+8nG3KSXpg
F5YFFWhSA5g53Lu4jtgsSnO3+Mj5uVyRSio0cY1Fv9tXgB7bCGwCWy8dEp2OKjmapdEZ8CjY7N2m
7h4n8TJrHKi8Em7u9Asy8Kx+659TRxTyLCezEgZAy3Nwxps8/G8cvlfQCvQ42OrDY471qXy3PDbv
+vfW33h2kGaSAX1h3+zbt/+3eBichHpdDciqBmBWT/c4Ycw8Nk2IoktzPSKJaEkXHeFi/GlVcOGn
R7n1xewaEbziLp2zLzhnnd9e4wHrq+i3IIcwCgv6QNiqdBM4cL0Mps83Q4vK+eIONsuCDxvq3aph
JFFZQs7lmGmtP1ah6zptCy2/WGaAVHM7k8NNbS0rARUXIWbMkcftZL/0hOaYGWs9/2u5/X4AC7/m
GLSpecS27nn0zoUoXgB5x4Cr45+qfH+Yr9gWuuQgHbBnrL6i8rlhL2cYDpW4V4ovGMH6p0K0M9Ls
Ab3U/hx8nCzOhHW+v3pBDD7mKVJ/YsF5c7Q0pyXkLeA1r/SBm0EfnQMTDaiq2+CMjN0B6FPn5GS2
bFqxchH/w9pjVpouAcK9y+1ZTsgssYTRkBcS4aZho2dqcsZsTK+EsQGlFtEUQ+uWEKWstmcdVa4H
Uofm+rKAKTGKhFIwiPwcPzo2uADV5zz+Atr9TaFlppySaZG4pCLRN/tCsmwW3tsN2UJ47dRsUdao
xrR4zkJFpGcpdweqjdrNCUqYfaF1TGFW+1ohWYPhPjF09b2C0+wJehX5LyL2eI/9+KHugU35BlRb
ULYWzzOb1wRSrLEVFqE9YGUbuFm1afGqj5KgCkCpW8EWNLE9dlTm/PO4REK6wtw8yuyi7tFw+ZvQ
xQj7CBHZoscAaQbTSpS2rYssiyRKCABv6Ed7HlVxIcxevCGcHCFxbP6oDZYNAPGKbjpjvxqvUiPf
jXawUdXbTTYsWVrTDMnuM06m2fGY0Y5C3mA2KivjxLSB+13d4Gu5vz/eOtmU4WGI5X6Ft2gzV2Bw
OSbitysgBb/Ulo4WvrrsJO2vcWKtfVLYu1X8G5yBXiknCYqWlqsds0LyQ1g/7JpA4Yl3lkgekY35
7iefl0+5btG3xCUEqnQzSUQYOMAidEdjJtGgOt1iPbYEMZ+9ezRAhtyW14Qnj4FspH475vDXawdb
WeIQD8yiP+7q0Pn5iuiliHctNkSB4Cc+WdH7iV83zzVXjzqzTTpS+NziyId3zb+/mV0Ph0hAOPu6
JQimu0fdr7XwryPJU41qiLwyOxpg5jdZTFmI+EcAKMawQ8EeveO2FHkj1lYda8VejhE8iKvLpe3a
yjs3XSL1GMQL2/kgYf1SGAY5QveymnkYWqzTB+guegGbUYyKkUIgoWypQSkSwx1pVVqH5mOmyTi4
fFbmnDcxcmLC0MmHCIJkbtpy7lylEs6KB+pYKLW442/yKOXUKMeeGRVMERdCpSjp/w7Q9w0b6l5B
sOMINQZgKXOHmfKz/48lqp9bZwRp8mIHfR4IycnOhxyotqPs58ftQiJogv63Qs/mfPNxv5ysN2mr
ypsFVFq5v5JKy3/dyjeaJnkn22JnJFCGZu5EPLh7Oc3rEdq//nOVQGUfodhUe9yLwCnWDW97mYB4
zWetl8qe1qzs7yR98t3zDsY7J+kci0wO89GVsRnjcNUViIyBC6IeFBA9TUyTjn2O3IpnK/nCv5wt
PSyHMw6zxkmuErQa7tVGSpleapJ0dM/u8yOvzeDYD2OpncI1q358A/kRVcHMSIuo2vXPUGNV971O
G0LN4s4qGiW+IqjnlUXbb7NKASKOPsQv9BQn6OWmSQgHBX1oobRd8pZFIoh1rJEW9hs7BtEw7d/a
cOQebdU89/kH0dk3sf4nFhwt7Ecq9DKNCk30HinO8P/tHkd2QZ6TdVka5soJYpax43OxMHuIkbnw
BERxRN6mzGt637UUZf0RmMhtRF00NC6K20r+023Yy4IQCthvs4f98aR7SFtAaAe85/T8a0asqj4g
Y/BXlClsib7/fm6oj82vZSpuz4BkovXCYn+Kw7kezIlhvVYLbfU7CIkle/tUaW/s4UWZGSEgdEeN
o4sTKib9BU1zmP1woU+D86ljit8gMO97Q/kyo4CuJ9/llYktYJNaTNSJfDJG5faMw9aYcmShXJM9
d+HYsi7DMsIOeOwAQ8PfMcHMHmU3Y3Xkf2Gh3w0OGDP/MsEw04VReCT+ZvEjtdgY4Y0GP6gv8zy+
eiU4ubo9o21J3Cev33NJpFUxG7hFFqwRxKNW4fX6LtxoZYEolZPYiEZfk9vuroQmrr4dlTekLHQr
G2upqWND4qMuKZL0BInHQLkPQyLZMLaKtgoEaL3SIwd9BWeu4+NcJNJxKT5sYuGQAJnPYZU25EH3
I++Kml4nxl9o/WDelbG3KjM1m2tySjSFtYNNMlV9lfHQ4OL3W0A0dGAR2i56uRyHKqJAeXI4utYU
l3EHA1ATjmb0Oa+tI2WwOVwVoXHGM5QHwZJ6lrSOqd/NJc6A1Ltbvhoa51nrXUbN7C59k3qrGOqV
9xwuekmMf96f3mZOmgO81JfdvpcXlXxzFL7ddTTO8/tGj140tT5e5mFzdSeeMNaC6U/LlOVaHe77
WijYf30JCc1o+RfGvZ1h5I+J/K+UsuzKO14oby4KNKizq09il/1SxMzsoZWC1plJ6OXx5+AnvDfT
6h6fBTRotWOCuhsWHys8nmzfkjTnrc2E9niLnWw6aG49btLKVKldrEaGzkkBUTy6YixOASZ5TJWh
2g3uhr9TTqZYqHE+5j7UlJFYK+Z/TNLbBgC0o4kF04rhADx/CD/c0+R6N9reaQfoTXihTDE3rZVh
9lltGCgz0M8cPCLh42uCEILFcCRSIPmfd6pzwlaBlu7XnNTzNkAcCTCHk1Zfu9tC+3varHYEn7gP
U0cxehK2wmzRmnoB+VNP9BrniX4LuLGjz5LQGpUNhcyDDsuEui8RQ9XhlWrG1IeY8VDH2vbpuP23
DkDk8P0biwAF+mtoJZrln3NAvnWmJjBIUI2lHnBuXSlqbA4PPVSX3Cp3/T9T7sWZ171Pe9VKLfI7
RyIJjODJpTS9VYrOx4g3HigSEIhKxzalfRZIyLv7YORZO+JhZ5Xo2CbhaknmfgzmTv3Dxdc4bHCL
EVfvKEZefrfb4kIXmPjD/fP98RjT0J6ybtB4VBT1Qb0Uq1N7uy5xVopN8CEhEWVxLSKnXyQtnLpt
Ec0ZA0r7PubRafx268VVaMvyiwuRIdxK5K0JlvhBTgS3pUbaXiLewvYfgzMPbynCNr+ydfJI7Y4J
ik20nqZ/9iU6e5pC6v3ByZx+xRlY9koPHhTGPQ43vyTT+QqkqVPDDGishfFdXGyjnMAWQde27n4g
wNJVrFB9YV1fnfuggfqysyJ73WtZY7C5rCubXr3opPwzSxJr7vVD+n0rSd1EpJsSjmAvu/cxZZeH
2SZZVI9FQr3XXMpZrLqa3g004OeI8Dm03KA/Cit5G/1VeXFpcpoVQQvvTcOcFOOEjHRUfJzsmU+g
N7TEKbwe6A2xyLazMK9MFEMpC7DW/WA1a50vFJw2OkjSh93KIAndRwgR86kvhzeL+W+JzGyGZa5/
+bfgGntT7rTFXxu8kIBe1FLtC7XZYCVfKmfFp3CLgyk4dXRfRFh9H8XtPJR3kvFeElhFAop2p5E4
eP3436g4E8qA1g1Ol8IO2wpNv3BD7SJaU0lR/F7tOiu+FWAcRmCfLSK7ajCciQ18cXr6XBvzbMBr
7gzyfFuv9HGDQbZQSe1YP6nLLmH0vlY/LWpGCrJwfNxIlVDPL93ZM+JWBrOlmJ+20SsbYeQ+UQh/
8E5ujEfkX9xkrv10VOVc8mKkMLB5P8wkvTFtAwTAsE7IpWQpdYkti4Yz6AAY9y6NO75X5SG7tmOD
Ljn10YlCAH94mlFHPcqpfmU8w9oS9lET5Vj+QZI2dVoM2nAZ/4msweonPQi7oxCh6oKXiU3V3tTJ
zASbU/ODuG4AD4vdGk7mIe05is8eZ5junGVmaU24HB/ZtFoWSKP2VWIhTvV2kXQqvbukSAKKMjKo
FW7oIfVnkx0kMnHBj/m1Vd6GRBgSF4+EDTNF6LvvaU+ykwThgnHfkayITkrGgtCRdq4bLESyiTRy
tOH94hcVNqxRpTF3EgMSpuHSpnWKFivoO2kL6kOYNqBT9FHKZJ7HSOLYqcEFyJfzf0KErmvyto1p
dReqwbw1qLVcJwneGzUSoPKEtChDVjMnSMZQagOOFcO9nSRQWRii4WlKsUzy0a6DVZIZqS+LMuZC
IUfeGfB1KCUQEsTNvDUZzt0N/ZfmCvOUJ7VqDKJLfF8FlEJyk+ZDckAV4a1E+8jm8JR4dyILHPB3
G5RduOcipiTDtj//tsQ/wdI40Co7H5YiTfqYGiHAIgIstDdsFf086AJPsIGnXOHEi/b5z3igTog2
dBZxmpdFNbCRGoTmeJsLVCYYTIEltcpvRE2H6bT4lJMK1bgFOcvPcn3bPkCEVcDf6htmVkKj1eND
43BUWl0vRXrmK2VajhaTM6aJJ5mWp+0TNlheiGaiSfs2z2KvgZS/9ufBsBi29q/u9Tk+p9P0uQwU
p9WWTumh9slMfaIh71bHhlHyYv0JPML2NAU/pKuhdOxqBBA239QIvULs7choJoZ5w6faXPR/r3KP
pwnE5tGIWlk2So7pRlI8FbEdd7FexQiy5Fmevv3t0pEX4DPPfrsyw3syQxPh/OWdOwv4F9JfG9fU
xMqqFdsT0XoU9FmMQoDJOVqcr6WB9PXczlmGTjjtT26D/h01SHJ/vFk46Cu1NB7Hth5eUuhJKsdu
1VVribZ375PyK4qng1cKZQM0y+CRHhvrqmzpshC+T9Jw3a3x/RBYyTIRPyNi2wdboIZ/V2jOgMgp
NOgiTZWWiI7OpwyO0iNbYpti0kV+F/Xe7lbim0AokFim+5nr3Mf4pWyG+7jDO9kmfGZ3LjEYO8Hs
sEhMgHaG5Z5FPHKZ+CgzuTPZ2tgvar0Iu2bVTji4v9XYHAfC8BZ5KKJWiIA9rY7M+2AqKwqxnTMU
bvUsHkcJR5pJ4s3kvAeqcTjyRn90F3oVWjsVuS3Hxhb8vGJk4tcgQGSt2m7qDfasTvLjX9BtB+of
BugXAnnpdztMVc0XM+F1zG413+JXVcyNSg9Vx35AB2IxdaRTk2JCMDfwBqEmdDq6+qTi84NFEnKe
ZFalxpM5My+7r9/JowQmoAQPq0sbb9BpU5YukqPv/hlbwxKh7DKYyr+CzLRMJnq3owLNWLV2mK5J
96SgxEaUhRuvNqjjomSU53r7HI0/9E5LPSU5IOT+zBM1EhPqPwVb7A27YLU1114Tlk1ydgBrBun9
lAMS1NUJZX1Lqot6muInOIIEynNBui45ZNW1Xg/WJ4mbvKS0lftAJ4ZNcEXuSdaJLSfQ0CkNOJLk
KGeHcathYN2ESpFrzkNlvvSACTpWJ0joXPtDJb9KX4qIRDp/htNsg3atkUIgUQu0ayJnGjB+vO8M
+VI9H+yd6jfFiO7DKbaSVh8ygFbnTr+fpSPF9FP+wCB28Z5RwDD+xRKoqtuL9MBQVTX8ay4EYkO1
NuyY+TjRf8OXmZq8vRrvd6Q/PLJUyFwucA8ZmraLpdnHsWLngqNXGAZXqwxUbjtwWhfTJuMKJYJb
dslW0RMJLsdudakdRbRQ98cRoG5S/YqbhetDAUcFfI+lOrozI6UfZUH+uxJZrotGnYbD7oBKyK91
viEVeWzUPJCr4PNMGgnAxNN/mlfeYzVayrdagK/heXqhIZLLaKXrQVrrnFJmYrCAFTxjGN82Rwg3
nyDChauPkw7Esssy93Rio9I+GlDdVNXXXYma+V8OkCtz6V1V7imVKoJYuXk+k0SO3OZUOUwVJwP+
Eit6QX5fvvD5k0AzQtjOlMrbLW9Endmo1ovCOx7txhvQjp5mA33CbyZ3KVbuQUlXtrSLikGExtUU
zWqMRFbhE87Ltv27z0k8iB8dxfxbGOUHt8SgFpch39JoQp4n07eB1SAzFTyRehWeLsprKxBLLiNB
oDGpz9zddBvpFZ4KpJ9exZcisjNkemIu9213f3vBLPBZjkwE+C399p2b/P667UNepP8XcfnVuk5V
u1zeE0B+C36WXBFGyIFMowqwKR4M/2ih8qIQf7ocxQcPnazETCp+agaY97RToCW2UmS9hPUmV5ne
MbJdLONCM7JxjcFbUayI/Wp5Pi/4oJhDtXP8WjgBQlGRnJiZ9LvNAT2oIC5HDZAjFzW3frFIv/Rc
5Ic5/EyPPywyv8zNTXs8JI+0NnqIhoOSuLNJA97Wt0PyTQVC7C2n+1nWBHIti2sG/r6rKpkuS1WN
nUgHprghOHzKSx6b8p1Y4koM+qT8RXTFVCbfgdbAzL/mWvHDHJtmet0xzv4QD2a+PQnp456wLgc4
x8Wtvnk63wjE9+goh49w0Ze8yNOe6fye/1OJhZJabxwItntkrn10DkCscrcecxWXC00I6JDY+tjB
vBMjvwXYxCdlshKuvPcLAeQSKDV7Q8w97183pxbXrwMbm5pSfvbAO3NnfOpDaOJ4uFq1koYUpbXq
a1uA/eoCVXAfHyB7xmMTTvQcOWYOSjZSdWWc5FsbYDuRbq7AOIsQ8SYkim3sEm0S+c9g8ztV8RVP
fx2YP22eaQxRlO8a8EeMzJBQFQB585SoMTDcpeutK+G8yPXNHYNSCUF6nH8JphFw7fpig1lynGsz
xhsbXde8eHV3QEBg6jsOccF4WYLXAyl50bV64TXlr5Cytnm9qWbsv/FhkuAk4EvBEM8dildvUNZK
wbCCXi2c3eF0GZUBXa4k3bD5HcoxRsrKBdzSZPZ/TGdI9jCEfPsJs/mXTcgLsmgyQuSyu+Szb2dC
KY3h3PM2LtEfdw8721GNW/Q8rUjLnIe+DcxYKzLNN+YVkhvIsh3BB2neNBs0JL9C03oBeS4WhkA4
A/xsNGsoRrDofhVwAeNEN7kt/p7W5rn887QbeiE6Ogp77kzT5jwln6XdKw2bQhGuFGpWFixk/LiO
/06iBr2Kx+iy6R+YvmDKCL0MJjxzGflVFPvzEiq//puqyY8ZnvPkcqot8v5A5/hZtQ8FGM1uqQS6
6L8QAefAQvILdnCqrLUefVv6QWRdjuHcAxVeE0tgU/Mr7w0Of4dVLr0tCsBgPluU5P8PRvI4Is+5
oD84hSBsAghi9+WjOysH4APS5OPQzmmDbo7ENF7t/TvSZ7G05NVDeI0jcbpGdA0CeyFlSQ42qvq8
ah8XpLsMAYA+CerpZigwpD3rDiwHrfubNc4XycMn+FG8kwS53cKaMkyE/JrgVwryK2L32jKUtyiM
6oBsmWMAYi0OPwm9JYxSWrW+lzVnDz33pCqPN7AAXkcWyHk63RiZjfDb3ghasFgcMqhsMNRUHEC5
H00hBtJ9EXoLqwxO/6pSbH5eZ4O1x/wWUJxapaF05/T+L2WfH1p2frqUbe4MfoATOYULtEenahRv
/dwCWmIEosbVPZnvfHJz5shc0dzS3bLTIOJ1TXS+BK1kA09myB72oqjQXg1mynhSq7tGNPviXDqY
CVVwFj+PsavfNE+BNdfFSzGnHGI3UR2AZRzbX7GPd/9Dmnxy6VTDxMfmKa5Ny1HXA6Sbh39ZiYKv
K0VBr+Y5kH0RiBKOhz+8lWSkDQZ0K44iroAuSQqWK9+p3H7SPmq5U845MyAD4Y0RtQNOLfxfa9ji
dkyTP7OrMbyPlfxIqDh8z8yNU5kw4Pb6CC3jpa9sjl/M8vf1tUtXNoa/bH1DxUe9QVGs7VXkqhC0
UDKRjkaHJutrqt58Iy3+utBLwN4tJlh9/fY5M66ajJnTwhfcYCbxEzwduvhyudXL7WtgJkHBmVjX
gjfSzUeFbuTFGBvEcZRQuuoFCJ1CGpHwXdStobjSFbN0c638GG89oWJy+CWpM3nEDnlekeuZM7mv
xEv0lujcdtdxYnjc24igCKDZa2KHV6+GKrtp+SGWcGOrtwe8c+kjcdurcqt3iU2JwVGNU/N+Mnxm
hLySPqABRNp6AI4/DTL1cw1sXmb1K77h99v0XaHXA9f0BHFCTFRdc7HWyH3spcy7VAKlq2KDswLE
7NjtkoIRB/SRsHeKmldkbrBeaK0YhiFRbM+US4vYQkl7C57fJG2LD0m11tuR07u/mjmF0PtnqVvA
SVaazycwQ9G3tVeEkVZHV0ZxXuFWcGBO06AXS/eCpyGc8TGbH/mG2ij8gdFRAk/GXaW2BYnSoApm
bl8Cz6zl0ZXHvCxqYFFisyoiuw805op56uPOxGJBe0jWSbwUk61xL6e3fP8XLIXoIIJwTnpAGIJE
vzs7HDdjCtPILfI6H0A+j+rJE/w3x+jyuOTxgJxAaKOdq40DudJPgSNuTC44FsfTGtPE2sWJvaqA
dZO+d+OuEl3T7D6CdU/YaMSG5lImEp/ZjxU2FwQpe4KA36WbqAGVfT911opYv2RRO7X9MiKExslt
UktDI3feUMqNZDXvCG6/urX5jmC3JDpe2dzAk7I1oVjht8ed0QqQnz/BYBpWnZE431Hi3tFlEQL1
uMyMAiT0xaMsnU+GolWOqltpEOZAFZ4eD2CV1/8IsOOPUpmk/Q1wfm9W5PDu63gZ4mXe7AhLvBnc
DZ0NuBXi1rEtrpF6uDnaBuW8bBSyU96UMtmH+AsymMVCFAq63NoZrNcRuLc/VfTOEPPNxDp3TqEh
RWS03F91kl+571ACKluYNzwAUHtM7AN+aOLvpnpjF+SCFU3PQF5OK1gpjoDipvNmwuU99mowdD3b
7VvBttXJ7sl5v+qaPfuIJnNCHzO/iyap5Si69gGklOmaHGI4nnuAiNAMMqLKm2D3zZnnGTNL8XyN
l+HEmca3flV7/fOfnZUT2h8tv7r2KSFcIOfhuLZ+MtXVHmAAKOYsf+P6gwc4k+3iAg/qbBy0lFBG
KKgHQBkQP4igOlBFfOd0r0r+pT8EFWURf3bkS+PhbAs2fp8D7nsF704YhWvvkqmpIsykrED3kRls
4HM4jRfbGX/Fewwfte8S6E05bFSYIEUQCMFSPBsXepO3LgAJFvg6FxJ6n/WyeescNBfEYWQRC61a
e/8W2PU+0xoX2fobdVtISj4Inyf/gRXIfJT9oz/0CXbxXLCyP+X2Q/SGEhfjFcWsDLS1kaPOx+aD
ICpNBgY2BkSMYxPomKkjuQSYFH8ypdNE2aiRuBNHHhanpCffTZdnCnlqpB7a7MRU+aVQYLp1hqo+
7oXwThL0e4T3Wp4MJJRiVLsvPtZr1YBxlleYfygk5vxg/sjSN4NSc5PYzQADCLrXD2QkdMZ1El7I
nyadvbsFKrAY+zPd477gtcE2R7vT9KxnhaTn6iTNcnqMGTGrv3Rt+QgN2nYeVBYtZDuTDDUOP306
VFjddcUEdMzxL4b6RmJY4cTUhQFEmnJPm4W3WmXMpUu4q5BCL9iaR28Tk8CRkYTCd+WpqR5Daals
eeplVY2IK70vjMbuzaQLvuMzJC4RUL3UAaovre7MIYITd2/YINyZdgKaU/ZxldI2hvO3rFR5n1LS
fikPk2TuKtf0/Pyfgjl+mKiL5GqYEctOVqFdInQMpFjbKfG4kXoBrtmBHIuU+PLjO1BVDWyrQ3E5
m2T1jAAjhY29QoMgU41uc7lQzXf22mugEneMOpJpKXnvlqzips3Q9hCOXYeNblvRc2wnIKUuCeAp
LPOmMtu+6sTsWQI7uay9Ws6Kk4ZhuNeJLaojVl+VhIeU2bhV9jRZmy6tFdvbT1Jv4Y79fDbJod7V
O1ti5ZGDtBrYUbCXO9avjR59+d0eXK0jESpW3V+RVDiOowfWwfRHR8aL2K1OFFGDqfUWNb0qT5bt
t2FHjzEcjOX2GKNyG8oQ3472nI2Gu17wB+vjt0vDoRI8wXNSFLMkTNP8Ak4UGwX1LacH9J7TAfBH
SNMCILBUvtioRBDSwMx//QCE76bolJsgICZcJfuSwlj1E+vsmkXD9ZWeG4dDAny/DKdDnUb+dJvw
wO1u3tvNJJIe11eTD7R4v8J9F8SAiDTvE8QEauTG/ziRnm8leqwyxbrTaP9t+mJqclocm0MnRdrg
wAM7gljQSB54Rao/qkO8eUiqgQvrLZ9vzsekYPqn8t6CGhsighqMn99VBXb12a4/7CaWUxcuZmSz
seriWIWrt/auB0AVjYvSFBt7jKj8i9uqC6KDODhw8TGqYye9Y2vrxBq1m+0OHV8x+8rS0o68Snnc
QtSA5oig/Yy5jbqfQ/aS4GI2ER+s2rfiVM+KqRkRn+kXWkDcjoSRJza41o/nLXImBcYDXUXNtbNH
tYjmSSIK0LvLz9s+2yFWHYPVKZcuyuQJwhZt8JfN2OHcxaK34pEp/JQuyDXAbIpsdVOw5fGY6B5Q
l7hkvzZLLlzodHU39clKYcsnBXF1fRQ8VCkVokm2Mqog7vd3J7qmMgQx4KqCsJNoXtkgSx0H5e2i
8RCk2sVeXXp1eHJj6C+lEqG3mLT5wGXT8oaE9Xiis3QL1MhH7RI6eTtqLoLMFT8WT4Ld7xigRrDR
4KqxuPzmtVsFt2s0OzTH+7uqroGhDaq+RK4udFwxRisAa7pepClyfJ8MEoTLvu0KKoiGkHnAyTTK
Uk973+PszpMxXHs7/fB8NxETyVM//c2sxe3dE4Gkm6SqRuJUkbPfOjwRlXSGAF3SUF/Y/YxwRoTJ
6r/gtNKCoOEZVDFA9xsoP2SS4j3tXE+ayrMzZajU3jF+8he6wVE3+DlH5EJO2ADjcf2d4L7ZlVfh
5UYrUpUjwPi8mSSgfGJEayHZfJPBaJr/fZjhnMKyhbmXUrWLCtMrIqDOE3ByPWQATINKl6cEN6HN
h98+tOosYnh5e0D3dsYgdrICWngvmr1ugSIFmLhLu79N9IM46vPeyAKAso/lTGxqVurMxjAUf2A4
RlTQAw98nkwuC6FxY/ev7mGOXlcJb5QrOc2VIDgq13oSnv2CEM7rWOrNe8ezLwm47rJIMIGodRSI
Sx87Z1H+ae4EvSGcxMPUaLLs8DUpKNIG/n8lBS2CGVtWg7sSac2+3Ec/Ph7S6LTISpMfBDIKqsIJ
+usnxx3vLVc7JhDEfdnQatfXCGUrNDHIAWoYHyMXQmR3wyfuXD/hW5WZnSYJDpWbbTlpTsL+WUfu
MZxOyRHLzYz/V1S/5+fvU76ScbOLLZAqiV3O+T7ApdNa02P7evi2IoF8UWfRMdAax4o3+lNbhjff
1RLB5EG3fckvDJxyTrYBQh0erpCgRYMFwyauVVASaVbh8lR+Lrft6+CF5sHty2LcL7lhPQHVwfTz
dLR6pgLuvZv10DNKDBdzIgb3ybrQAglflJebg8nHYpTsccU3+2IPUzXItowfJbzL5hwSruLDt0F0
J9odpbU4XDlJL9sBwjcogJeFumSAgEzDuCL6lSissrAqPYZiqzVZ8PJ4oh2m/pg0pazZJslitFzG
1MwYl4Ox/vISG+qROu3wIOngui0Cz3G+a4Owsqynl/CRzQCj9t/YiZZ9v9BTESPU13sXUOBhsfYt
YfOzgusDVK6l/JrPWNT+cq12ylaxOqK6pCxnS1Dejhc9yJAKyKRelkDdTwx005mrPpt8beyt9Sjt
aC3D4aNKutEZnVwaiGje2FqJWTnYIihlZcwIA8roiVxvNpzLwCeEgdflHlPA3ILfy8EmCPgfYILw
AhVKLO06P6AgPsSGEwsfTKbhSrEhxvTDIEiAocOcViyXCrWby8KWZLSTsh85i3QIl0UeESnYnSt7
VOIw3TAm6FSpCejtLCFRSu6syEw7iRDqEHo9a6o93/QlYJbmBSh9iqdxDjkpVGbdjTDAsLsRooWk
cTWHURY/jBk7K9m1uDorF4/DMVn6GbSKOcP3gCcZUkOCkrOpaNWwLvoERQqquLyy9uAYecOXZVM7
uKgsKR+yhVCQwxET9VvCeZiy2JLfLvZfLyKUW9nkkQUtqBL2sLGBBEAILCHUr59CKUTUF+mbBgnD
EpKufWrLAUwaRF23b9K9eCkdBHPWiLWcNnM3khXUEZohYcAmZKQ/1/wYVYBuEZFM/dNYei7mKvaL
UJ7LiSkQr4/Dz7avZC1WyFW4ZqOrdzdcTUSmqt4Ex2edDYLjT2jlmKhyCmOLSrVcV6R3sZ38BPiO
a3tMJnEPyYUHd35sbtNAF8tC9LXRwLWMZm8L5NdQdyN+7RC6RpNuFOKDaXtf4LRTQjRHxHE/EJfP
YQYi8Smf+sgH7ARoAvE6FMGE89u06oBItzuddJsR3b7qsNm6c/EOc1cqqSDVn8wdS6sgDsiE/zY8
ZBgiS/+a85VYf9/R6Xt+rgT6nAdYfZsiQ8yVxKwDbtOXHfhkqvtSo5HEDTV8TNcWTb4/XHndtDJs
jGLXvyU/gYU0iTjtBPIDzOiI8XCfmPkSNRz3MSsK/wL4DrF2z7xb/aTy/sPH6kzwFDdIYYaK6QgT
/PPMM3/Pfp45ca+K0wRS7ize0sXuFFNe7mRPhf38z99/bvt1NJ+MD03LD9DTnFI9aT30AS894oxH
inAt1omkN5IWYJ89Bhij2ou+IFyLj/VOltK4nksefHpaL2O3Tun+tCFKPrqkuyJj2ccAkYdlf/kC
7tDzHH3yvW/sMjH7HwQS48SyvbWBBqTdDBThjWKseUWUX6Zd12cMbyTHtva3eMmMfvSQKAxmc4bG
NW0S9wuI+L2IzJFZ+zGSoNnZ3OL4220rui7tfSISJlabrSzVYPsz0XX055DUXno10Koo+x1Qb7oO
4MX9D1rgBC1J42C5pkziSBaopEsK1EfZjrZHAgK5jNTLI65bQwTeVmbCF9T7zFXmXu1J/k+Ev6O0
Ap0M3CluK+6Z94y2p7zYoMat2PG9oKI9XMGrPZClI8v0ki8wbyxDuRZZItA7zu0MwnQGSHr5dGiU
EgUrs9eVzJ/VvJVhVdWvbLAx/vsXBhx+c/q6vWiYtVUWHMzijyctOd8tDp9CO3R0O575gGK++pHE
ZiC/iiTfZxJ7ad2EHkvE64LMMNN992KTycgoIPP8lEGm5ObtF6XAfbufi73/4l34Tk/p8cL0+CNJ
NqWtU/lsk0Bl7tLkSfFNn2EeeVfnNO5furhQ3gIM+OR8XzuTkL0A77n81CgCnEarALWN6rwr3Auy
YE0x9rBda3nERJHRl9Mom38D0qUYJhM4W/A7Eb651wmD8ybBH49Dp2gxBQtPYQjLxalWgqiuBFAj
UE5iX/DBhJ3jNx9XLVAFPw2V0iEQVYvAtXWtcYfPdbfErQkTjMwT9QoFS4vMUeWD1hRyVb3sW9Py
dmvSaYrkqf86/0XIx/f5DVSabGy+AF1BbBAQu77m+Fdbr4o7VCHFCj/Y+7Fq9APRNMOfifZ6WSaB
rfEw8oHEDsYjqrDjKA3D1CFlmgxvUUDBfIon5TyH0Z+ZvmZJBVzuP7SFlPrygDexjO7TxHChsVYe
S++URU9O/qZ2QhPJyDYJ0dUbymliyrayeZtAs0K/bE1hNQuBGZK3YRJ1y1+p5R3Ih3D83zyD4JxB
DyKyH5NmZj3WcIl0kE5GHsQa+YdrdePOrUvB3ePZo0CHba6fhrG4haI/HeTayD7DYG3QpDWKrioT
MgTSfwv3pRsXqssa0roISceYm0W1ahqRJwrMKEPdF7EmLJXPUu5u6ZOHYZbjs/BW5zpWO1wEfTXs
wokf6BzpSCGUagKPCuVGMDgBTz0BzYNrsamBAg0pGUSLyD4TCbkI3iQekVoAHo5SCUqI7nm5Eotz
X9Z8ESpi3OJ/8TkqSXD6iIDd7RvEwfxWPaVWEIQklcyzcOkwEMQlL1OvWG36tE50CQQFV/CnzYm/
lMqoHNdbUdKASNPa77NvrHS8d1XllxhuUXuK54WjNRHUpLfQBx/pxp3L0giuRpiywrY+GC5JpX4F
rJsziqnWAALaqhika/E7RTP7fpgBDAT7k5hbMoBDZCBlYcNjQ7/Z8tY3C1Lhbo2358M9uk23Fg7j
xVo9M39T1DDiTLnZ6n62zPKhFnK1ihAROXVQI6oBsGoOwty6MOCmU2I+qtIGX3ECq5oNLb1mzHy2
4dU8+dg/WhScmfISh+HjZ1QclpC3bG0kykZb2QR9GMsJKBpoegiZun/si95wdGg7hlNMsgMcn+ct
EZXis7CgmZjjP7wzVJwlU6JHW+Y/fmkmlYJW0I6N4ttIwan/Z4dX7gt0LXhHigC/8BIaP4eiZGev
1fZ09/YJ5V0iPUHUBSGs2cpMEXR8DYjJUi3EUeAdJsp4kPnTIO0g1cQETcBTdqN/3UMWq0mmo1Dm
/kiBL+8HC9/mevyaMoV+UvsQ0cl2SrgeeWIvh76blT2/9FeQQhB1p88hCawsnLNSV4P+9Vi7ylyZ
wzwZ2UvmgedngDgmH3ovL9pD+/ee5ZKaWR5Cv/Sufgjtp0eCVsSCKAPbHQwm6UlEoV2sgdLNBlNo
7sWq+5gJ5v4bz3VTuuUpcP6ZuCPOk/Li0kTdslnegP3a+UaW0Wvd+j6MEN5HwFPoz7fRRD0dg8mU
TwI6NR7OA83v7vj9gNeRQ6sScRxPV8LgUwnoiK1QnPfdb2T2zwEwBZDr+Q384loOQ+U4SzBHgFyq
+ucjnn0q/HgKLesCIk8BO6q8lcB0TBBZlYkyKS/TeIHNPgos9GUQf6Wo0lCNKaurlfWbS8fxW3j+
41ZuMm2CToP7vbef3XJ3i9WA0TrYbdflJlL4k+xxWG3FGk0SEnslBOioJG6lxWSH2HYQVrGO2Rq/
Je+KhigeojdGOc1KGTOxiIOoY5rV4NCZ0dM3xmIB7TtbshLlNuCeqTy5Jaolgu9yJVn1Ux5HJE/N
xAdOfZdpkdZHr9wsZQW0HFNyiY0BiwPbv+FBP0YiCbeYpcjlGMFVpMHDZTAzaDTdrdnsvG6Ex4O2
l4fJIfihEq3H+LI/kn/ulmD8qA989qTf92dFdZhdxgu6PmdS3MIVjW0P2zFF04BHv6OigGv7jLAb
tDUB+8nu4Y2V9+J0vXFxdz4UpELWPuV+YimWBMEm+3ZF9MphFms2mjuru+XDSGF0/A3Elmo9o0uf
8DD/6s2NfP79cEL1ZZIKOnzyfcj7JaFX06l4DDrIFe1fJlcpaBeQu3pWhjTRKYxbYPdNeJm6hHG1
C4CNmoM7PVDZfFqxG8lBDHZlNlHJU0AG1SJtm4R0WVcEyMOjoR8PVf+IZjouwH3Nsb//iwQCK7Yc
a51S2BBRU+IVQvWThmFKYC6gFiKb4tuFuPEywASfJHxd55S9VY4Zgb8mrh2bztZtl2mlPH/0gBbt
jOePZwvS9yM0CrVWMZxdDM5D0LV6bwQa2rvBAYxR03lyMnM9+cQKK/m0QSC+CN7vNyF0kWDMLjMv
NwQNiot+9Jfiu5fkw4SMsw+6X4Xei2tAKq7a3NjYehZozwDoW0Vpo3GhNJ1468ywAXL2M3RanRWx
VlH6EldDZcMxWGaQ8s/xZnmZXMV7rbhzehQ85+9a8oa3SaxBcDZeSBsFJTvhvFftP2zIXnEUxzAp
KlUIp4j7OR/+qFD975ZcJF0KCRccTMQPfwOe1ZuFteG7ecEBKrw8Do5ntzDOWeQMWXKZDitN8sRL
bVCCIlDyr66iXlCWLyEYg0+F/TKYw+JesyTt9CuFXr5oYYuH8c2Itm2IixZUMPU6FUMp9KzIgArw
LifeWCZcEgzrUWDhgAicDeilolH9a7vcOASDBwFk2XXcbvSs8nunIifEdXJlDQOLH5tg2H/SiONB
AEqscUZk/tLvqMEaSXNtXZBeRw7zYNqVytzyBpFtsBUDhKdGzJjU7nJY3L21ZqE4cIo2uXco1Sif
D6aDmfgIhoJ+ozIyE19FtAeN8XudG5adM44H5u53c04eZ95ACNcBg+M4o6yag5DbExq2l6Bfwzm9
JcH3WiYqwwYsj4wt4hinlSmGWSq/gCa/AmNaClRSmPXb6NiFEf/vXMUEXj0JUHtxUHqCQfq+eQcB
0WUz+tihvpV91Xq6P1yyc3ZYRmB5FA5H71Sj5bmE5doP/y6cZFsAke+tFWSBxmdhefBYSj7eoVKT
N0Q7l5a9djX7jjOqVpi4Rm4lN9AJh+KFi6YZu0R5b6v2V3CMK0lN8DUEIJHnJPN6mnGgbfLO+ISf
DrhNwhsBgPkPcWzKq3rXcdtE2qeLT0oEMGf6LnypWZU53tRrVFy20wh4By47VD6gKEVf6XVXT+dh
eMpzL6DdhN7LWY7tsHqIxqDd6KF0Ty+hA19UQwd4jvF65RuYT6ih24PfRbnI2YgNsqG/aQiJxam1
6K28gBHnXng6XRoSyC97tp/enZBMz36djz7ELpWKqhrOiDKg7z/Z3x51y1PtLtUVn6Gl/fciGui2
2eKhIJNHUks3M5oFR1Mw1YzQlw0iANx70UPnQOxgQqXdRmz1NJ/Ps/k5rfaH/7KoTtjJoce22hOS
SgqktL5gLpCGwCFCEiR81Tn5kXmjowAU/8JP9cKVS81OdjeXEwp3/zUCqlg/VH0eLuVT8Ieodq+Y
kOgv3iACBricSpS2x05q4lsdtjF4DNKbWH12SpbUKlTxdJWveVjbXscGtb9a85XbYno9oOJVl1T0
MTZOJtN9TR+UeVSL1MlAcCVkn5J1dPbDh07fDC5ctTx0/xGRsYZinaRv9os3OxHr9nULATSYntLu
Lczh+nfLEX1UFwBITrhHqXkYbAqEiz63dQOabsWiP4a7fwU/p+AShaR/B6O4q5gCcaMy3MRkVxek
oJ2UKLEJK7ZjPKIZnC9as6aP0ZwST5kNO5mdCJ+8+mcvsLysjVeDnWtFzm5mm4Se1lD5VMjkYqVT
yCXo4WgIHlF+PikDLA+GENMbqDgNs8eC3CWxIiyOM4hG1B2FDT/2E8r40EN6TqtgsbqZ9W3UTOs4
z2vJTd15q+pRCiEs9KOoAYxihYiuTCaYA567Y9uQgMZnEeGQX2ycHggu2xVNIVb8saH7QWJ1Our+
5CMCg9uUCJY503vzsGMmeu5ohy7CGW1hp2B/4annjmY9HyVBxasZAVCYLrsyA8CimzsZx5u/YMRS
xz/LEOaog4JSr5X/bdAky03XWPfvkmCOgUWo39FggkwgviuAnC5iYwRKvivpRxRIX9qoTU6CvT7E
FV191hJSDGL0iLCGwhfFc4RF0vm8/vrtv0Jh8V8lG0P8WUqcehNxSssfkmJ1I6e59lmBIQ7MAu5t
nY0C2NUtr6+oH4y15TtDAJI1l3yZ83URBAaomYHgyXJ45BVV4g/tkxKE5qOtFSf0KOI8qxdr0MHm
b08qN01Y+t3TvojjO7TCAPrYsW7mUaRrC2lDKVcezXGlceTkqNjUxbYkLcsJzlcVMhuST6Wx9FgP
4blcjq+xf/B1M40LVHqMnsxjqac+fTqP7n5PWkFYLsxu9kRssxZFZaxMxgrm+tWKpi3bvw0GKkGl
O6Z1LSp/zUN9vpVrfNEUcmP1z4R/JK3d8fFfngMs3I8QPAQTCTMVJa3VFOTnnObDOhYoKMkhYlQu
C7YUxoFNMVLeIaHLlx/DPJ6ESqcrotGqBVDtnYGqhjgdW+SQPnASbucAG5VgzggKGLh/atvy89Gg
MlBvM12sX2sI58xQHAtuqKZ41fXVhqCMid4eqrhEYRhlKwfFZ78MeuGywMRXL7BBC3VqOBbtNu1P
r3UjFuBwC1wp+jehBD2kVYcAvcFvE+dNQRF6Z0bynmncArfhARO8sUHas0w5Q6fXIq0vkSyVWvXF
5mJbh5JkuPVpEt2rNH0UfEpFgw8Mr7itkzGHCn9Z+EIWzyGVr7zcjZS6urq5AsNZugWlQXr0W4EL
GSZIAF9hAEt9hj5zOi6+85h35N3QKX7x6M51qVXJyVBADXS1EAgOu5PAfWOt1IM9r/eVNmHXTEz7
pU5qEAPO2mm86flFCvB9IqbdN3SY4D8D9ZZcxx2ogYi2PpRbGWNn9Sm9ioTUse1t2YBWkFysYIXh
bNY/2/HfINinx3TCXLZCHkz6dWdRVFRcDUOYTNSrSBgS53f4G9GrTnD4BTPO9OoTxm4KemHiQhYt
R2DY+CLxQrn00bADHiTiOA7T+x1TUNdKm3/fa+SFamXgo2VUWV2OWmifSwnLk4ywDyUIcbwwqskr
fzCvdDZuRCKNROHPkuPYgx66cQBjJmdqbIySFnLKCi6+jdmk6j+uFiFicejfHafU3TqsFCXpXddq
67g9Lx/bFGsULcABQ8nDQOOlC+fsWaK/Xy/zHtOZ76TtfdYFtm/FMsSAtpeHzle4rMKq9x8cb/Jm
VEFU17W7OueaEibqAa7U406nHzAx5t6C+Wr7zDWnIgtDok7l2yJFQ7A5UfzXuiBdnpcd4XgNVLhB
xraKjZy8x/TKwyphAKNV/t4lRImr+61kLXM9Oghu7DugNp42dO8oTLwD3Nk0vO8vavoxZ0RQGac9
bkQrfpZ2mk0WTjQ1xSqPiuDtr/v7aev5fn+NMQZbKhql/Q8+xJ9LYD+FvCF42fFpRcXrZzvBrF9d
XY8Z7yOLpZz2eh7TSuoMnxIl/mcTbjRV8/e3NeDQs8+NS+JR3meWZIj5TRs7IKZNEIn2+pEaYRsd
lgJPlsixWe/f0zGSO0LCqjU3rmbhSFgfsObH+Fyc2rpGm5zw4xI62/4Xfd6EcmcmmZ4nmoOfzIX0
nEJDYz+4W/5/LS4zjnTUow/dCeG9xi/g2dkU1+M6jZMpL/PCD59H7FFVgFWOPM/r542atJ/g1ywb
WLxtnQSlAA0nU0NdbSadFwVRNHzh3/hV6oQTltq3NQcnxGsMoSTZyT/seSwTbExhmUxWpJTIypS2
MCuV6vziRUU7AWfzeYBFR0pIB6DVMVC0qCy1sRUfOqoJCOP7OsFZwkOq8fDAHJ5jSfZfhiBoWWby
H02RKZw8RZ0R6EafKX355trkxYq9JHBt8RjSinwj+m4az7vyCBuAqIhUdO4g6yyb53OFcvD0VoCO
8McOYmkZR/5jF7nO6Che0zZv0/8bEzVNJqeHDh4mq0s/lYYPb4HDfi8XBgT30NFQ1sA/0zouju2J
yT5NcIuQyPyhrppYycSPlzvA/FJf5utqBIWeEmNScVQ4SNkacVq7+MWBVUgvnhmRvvjRXCmP9CYO
DJxVypCy5OOefoLpx51ZM4PDRa4+T7ECgwS8Zrqy6V6Wcs3rOlIzfjgb2BexCGMyYfV1/ENmm62c
S8KAqx8fEQ5/l4vUgYB8Bib7wF5spWYi/4AJfEkl65Lc5qRrWl7XIXuByAs2djlGFWg30Nlb+L+L
ZWymQZ0sBScbQc9Kcqi46qNqeEF8flTbV7xubUe7f/nxT7BDcvBDqiW3i+JorUs0aGQzV7nhxvZM
3kCr2sglWrPEteLFiQsjuAmcnJd8lh29bC25KqRax8+AWsz1DRsjD9HZvdHKmhrdygVvyzypP0Lu
Ha4Ry5vY7frebzGR4kkni4ziPBRm9qfiznyTEidaFlJ9iKbBttAYveZaQ44ETQSQVCpwCo960nJx
3+Y6x3pspG+6j9WnfWw4gAkX7py3ZakZAVMpmaqgY2wdfAPXyQ5YAU/ymp9qUKD/o1NphQEyBHcy
G/293Pab5faBETRXFbaEJeq4esKIuqCbW8eHNUVNGFW9CKOjB/zZvQ3P/dmGhnmlBoNruLCZy1On
4C8Djla+boysrJ+JC3jrJ7e4nP6L7yrLuzUa+CX2hO2WPefX9bEqTp8NNl0+5MKTBCtOrCxWhGYI
Y1n5zpgv+lPk33qkZJo4rVfM3yy6FThSNAdZuMyzjU9NLnwgI4J4LF7wfs+RWDhmt8g9jV0UbJef
ZuskkmFeNCUe2cWK2YwMW2QP4M6wQoTtkFD8vLX2Y5JCwYVUxCtOTZLxxX7q4c4t/vBjU1/iWIbN
bY6G1S5OtM9g3ZZWFHJtIHPgl88NYHUNCVZu4zHgdi4aS/V0eWY02X7kQxf5U+ZTUFVF+flI/kZR
4voKK6Xp7zLJiFYa0HZTK4ocd/HomSVdtx5zkRvuMlh1lBuC3pGlvStuvLmRk+4CtVLDZBpJx3us
tFPxkLiqfSam1BDLOKlCjdMSCZjIHSZDq9wYDKOfhGEHOho0gVi0dBA94ab6BC8lvXQMPyvnnZn6
oGb7h8zh8yRA1IiH0IoiivHROyxMZhkyuA7hOS1sQAHkeD5En2cMl7phtNvKYOXoBgFPBtITdj4D
t9ZQfcL/tv0NkODuih+1HjiV+7L7wck0Qak+JV8BHOJ8f1IGT3XimZb/LvB/gDSjRrZ6lVGAJjsi
Fp+toT83ZFh2q53Tf/rCqozBPU9lsmcP4BDqztQJeA+TVKRPusrEs4/yMeGoAJ07WQ60D1dgW5XF
6UobM0g0H1fzTELdlBGRQVCxY8MSe0ijD4Iub1QnaOvXxaS7NeUKKUjOaFGpJQqjaLqVK6rhNkqH
xblH84iqLPn1lC29j8ocB6Xy8/hOyHZKf+dCW0GzTqSBoM/inQEdLlMMklXvN6ynjVsMUED3l6Dt
gFpUj0Z9yAXtqdfLw6gLyLkmsZ5vCsQNRV+D+oPSiSGU2JPyQDsUGUtwkNz6/jVDJHhPULTcxOiN
bhR3BAV5w9zzg/H6OiKZDAcTN2eElAQ9KQPIPGEvCJ3k8mi6QIzFM7RouaQNgcfRBMJ/S995+hHx
tFE1GP2TfD1jh9qIYo/ur+WfAEiMn58GjefyyV+G+RVFGpXxVdgcGh/rWoZzX3Xh7XjU699DsobT
/xKBzZyOvT9PbB1BAigSytMaGuD4s9XQ4ei0NedwuQl4KQAi5l4k/pz+71SuPhzP+QYg+6nOJ+2P
E8IMTydGaGc3Qx73rv2L2kPJNaSANsGWZxHbJ3G/ud6GdvedEeok85Y3stu+++fSxR3NWdkUoLUU
Pun9h4ph/RpYej3zkP0XyH8T5t+q7GrbH+vdJsJoeGeJbor3w1p5uKBN/9Br0AE3yZYGrwE/XH4C
snfaeIRALggQG9Inuae9U0dNRtS8eweaRUbzbTjNf/uQvaHDiJojk7gqxvdUcPY2iBpznoYEk79i
169t07NDSAk0rwBn+isC3aHrMhrt9NMmuHPMGh3nW8k0E0FUJY07d3gqB0Duii7E6G0peJl2VZWo
2NlQAm2Jp1bhTagTS5JpPH5XIWXtvcKzVIFzyjGZTNUsvnDxzopL3GVQeYihtdPFMJ8t5CX6bWv5
5Zhe8QBJ9sgZ2J7kl4ghYM/L6FUHmz9/7h6g1LIVSR+J+enjqmJnf/9LL3pcRNbmC5Yh41yyz+KQ
kkebEzWpgHNxEL9yn0ZsFjRqZMgFjHohuQ3mn+LvE+Fv0qXohJinV9xSH8U9+icnniR9Uf8FbCy7
5lyFhx7aZFmFaiMyxY6elDarBfhnhNxjELWzTpekVP/grPEdwNYNq77m6S1Z99mWtlF0aQsWHV/U
otiy3xzosjQw9/HwoPA2y25OaQLk3bYxCbZFluNzKVDSEZvPDfBGDDFfke9V7dcnz+LBLp5kVnfB
2xW9pztckQteFjxFtm5Dre9iocfq0iPWjYvH3kzNFZlIfHaujryMSB6uGndu7hmkTA9XjsPU9ZP/
nMgMJTMMfQ27zba+Rypj/pUC5Ivce3bqjVauLxSPRJebyTFeX7EenbXRNYXyxNt9Yf4ilX66ybEy
OjtQnZM7spmZW1erl+7OBcsp/bu1L3X55BCorP4BqC6nvwPprkqCHcKd0A0pGXnpBS4XLLHJjsxi
JLvbdpXw/YAhawqs+JG6ZzMM+GQOebrrrkz0n/7VVR5bzNVfLS8x3fStStskMKWcVA57aUu0z1UA
EfhpVONNSJOu54D04SAfgY8u0MpE2LgWDpSGcwj0nwkoNfqoOatDTLrag3B/05TS3AqRIO6fNhqM
hZPXo4GnBvjg7l6qufBTWrX05JS6fKs+hUvn6jQDUDdyuPoTcLFE9vS4C1nFYZTGFSC7TfQ9cBHY
Tdq9dQgDVgwUG6qJXvF8xjJbAJLlwoV0lCx1SSrXIHniXg+o4c5PKVm58puVzfnGTISWHux8/BgA
OO3xAAxNKDWbpdmZUeyScEizuSrSBafNTvlmoPULo7yLgizfVrVL3gycUKJR74to8OOhrVD/L++N
7L7MaeL0S5H+N76DOvj+GzKZ0sZOeIf3jQbHre9fvIkW1m2lwBUJgqEpOPigu9q+s2z4oVdj56CN
UTXSnJI0JomHkhrWt5FGNrRFkzXiRze6dOYyIw20nP/5NdoFu02/gyBLZSGJ71B/LbsfCjqLkppj
eVpyONDPFdvnBClFrzFIYSkDx7Zs1E1EmFPTOE9h92I3+5zuPOMeyaGL8owIkVxwppv8L7WmJ8di
m0y99E2vBkPx/gTAGfoXbpl3Y8TEidt7Q48L5LBdfCdR+9Lm+zK9l6XQCUgKDXi7ryTYuT6YRPRJ
wD3uO5+ybc6Q5bqfYqDddMVwhDY0voKKnILC3A+8M14g8mgmP3rlC5sziTOjHcnwtqosduD33RSd
Lum3sKSeuUL3fuhM7WSLwqYr/cOpMHoI8pAvy3oIQ0wAweCkLgToie0Lyosom5UcDVtZQuqc01Yx
rdpHM2FHbbTQ346tREdQZtoCAVe6FQtJILbRujf8TDUVqEhzhvqqeBKkZKgRupIvMMGABJX+A2EQ
MYWsXIN/o42T89JUBhXeFedHA5vqmKhjuQdClm7VgDs2Tp+GjLtv+zpaH5h41Nnem6DrgErb/yjo
WKnx1Sl5aXE9vpdzaG8/3wLQlFCyeI0mZXkgl9LSaxYGdv9MzOuhNxnQdBpBN1n5qnYD79KeQhI6
uMhWteWY3cElPiSvfPxGO4J0TTC+aGmMTNaoK8jv/eDDv8X0o4lQRObbn6yXNEQvjCHFhjSVG85h
h+qroDr4fK10n4hJpv7EfH5fM/okF0lnFeAYLD3HBF7CPxBX84m1KNm2jAAit+Gt5CUTDGnkysg1
+LNw7spsoGHVxs9cgb9+hQoFxbtPBIxX0mB/UuWrgEFy8AcIlEbhkx6RCOLrLMKscF0da8uRpBUw
HUnZDuuwBL+KtfZMR55guZIEAaxMCLX2Ofr4Ngb/DY/r+Z9gWXdgVt2aDCQ8VycVn5HMSefTU3/t
JH8Q+XqPLVV0AObFZ2PkEBJuo5W/KAl9FvaPJXtgagf64Ox2TZXv0Gfd9lxtprKMs7JOoHHSydYx
lWaQVl5VPwrf++zTt2U61SPTEdw/Rd5OYWBYUGZsyOqo8JMFH1uSJYqbikjygDSdoGRavy2mW9yv
sDtyjImileFlkAqe7mwJFcHG7zflgqmd5v7HXBBIijn458XA89NyF4BSKVwAI5z5ogBRLzwVWJsy
NTfw3cxmlZG989r/b3x24WsYYF9LW7h3XzQaoBOLpiBeH4yeCKS4MFz8WSzrLvFzuRDVn9FqITih
QHzpVjJSY3XIHnlTmbhbcRT+5aWW4mpysplEVaNDjRpGCJ+qjhAnBJhIFFkyWqUFe9bH5MbAxE2+
3iMONpz3ii0ifg1o707s7WuFPtOhTclVZD0xYge1vY9i7myXbm+whgOzeIXWHCnVQ5nf1HRaGkH/
lPMEgYYQubTscTGYu7dT7CwF32aW609w7pP60dA70/TcHOtm2sR5NaE8STxPbpu6BkdLxSBw0JT/
p3TJRaJ/SUpTYgZiJcnaxBe0UrEzkpudjfh53p1tpIagIS97zqQUPFRYk3c621uRfDtOXQT/DdXi
jB+YltsZdBxNZNbTvjDO49R8kQBtoxrU9h1XY61QPHhGn3ipSQoT+zPGZ5NngCNrY78OqK+STDZ0
ZlzpI6xcaKuaIot61wzs2+hGgNbt0T+utTMIRbOO77/272/2h/+EXQocD4nzGV+eomg6loA8rBIH
Zp42Rn6T7q0t5o+OcdrKYOXsJgmXTJvmbA+LH2EN8U9TPryio3ghy0XOtCSYIKwOZzVIkJHKMrct
17dCscevEOP/zKQrJnvm5mX0QANk8QJlu1Zt80ENrHh7nOtFw4AfR3G1TzxIyqpC4Fxt1EpQ/fPI
CL4x9/4RDQcbu0jr5QGvNqiMw6A3T6EpMyGVsftXIozXbwB979K5B8GCgBYKiuLpuvVuN99ryFYI
+Z5xIRD4SbwtxtPMZQjJzwHMZ4YNwIWQsQ5GT607ZBkFyd2ZkwogupV07cKNSzwcH+KWEjnI3X98
gW0lQLOVuvShHKwsNPKDotkedieie/wRvBJitQrDkFYYxdSWYTDcNKkwrW9qYPj33KD8ViyOHh4U
1D/461baFU6X9Ck6LVMU2YLUoDbrVahLmNr9ENWlp6WdPerQ3u70IM86cvmL4oC6YV4jqB+x8U2r
eG0ieUjGKsb5Fd+U4QKLBTUyCinXmIYR7IERLoElZcOCfUFH31GhKT7eN9AGwOTrEwcyMDH6/YkO
nfGeHWiDl9bf0nEwDIcc8ex/Q5E6NpccamnsOvk65UNlnT7COUraY36rKJZLxr9s353RA7XXtkVU
8FhkwhHcOF5jeTiENPpzSH70MvwVTVXEXoeHzGyodMHA0ty5g/0sWD/7E4/izMbdOo64+4MwQVv/
ZTOwsnwp0+1K2HaMWBjVLKdXo6M/7yemvzNS9RepQ/G3p3AXljsaTfFzVI5IrHfbuLmEwfhI3aD8
XbiPkOBSvbl94APd4HMKqm+PS+CMaZ1QZlbKrl2F3H4rFkdbekF5TTY2Fd500cbEwJi7jV4QE98H
nOfnPqdhI5l1Oh5jQW5CGO2I3gT9Y9/MdMm9d8zxNb5bGqy14F4I4dOe0gvEsjI5HUxGoWsvrJ+G
xayI27x+FHiF2FjKUeoxINxXOvMf5HS4W7Exk8n/6JalettxSQcQw8j72wck9euk6aai4/GDhe30
jQDyt6M+lL4I+rivVS++CdL7XW6bwkTO4lkbnT+aOBTmQs2i7FUEfWii7i5dE+IJuNBI1njlOJ6h
U2mSFGzdQjAGeIFlsqFs6ZKMvtnFC2POGt10+g8rF04QAP/Urmp2IQCbmCBFAiXLnMxLIXXfjc2+
UMewJrYPdSkfWxSt2+PNfhb5kJkq2lg0ddtfHeS0+/clW+Msrm001BPMT953dnjSnDQHr2ZEbMDU
wQ7gq92fhCiRHv0cFTBxZPY1S5gceyU5HDTf8+o8MSkhPJCjAQpzmLHqCTp9KxLXIl5++Ctz163t
jSxMxUOdcPFn06CJodRrwTQLlJrzyCSJ2zAtJtLDHAnQqdRw1od1R+a3Y80saOSVmlakHUxsK55W
u8KstemkqEw51NGoTU0Rups4drsQxkAE3rhY9nRmopgqXdcRmwGtl65m8a597YIyZqbKu2qLz+xA
FaypPVnmWEqUrY9rffnZiC4zyceZ8vrBQIuggJxzaGUcAvyU/fiKUJUs9oxwYKyzmrWufRB+xeGr
RRp6bUcRopJTbXma9FlMARIrtYW67NosoBocFCuvKsj3m6QLJmc1rxcMpVwLry3f7u22NQ+y3tN/
AhIEzdvP5IXGMsQEtynQyHsdhUX4OhUhQilDg2SLkIcL+JXS2df8NnJt1lv0VdHlfKqZ3o9Q8HNQ
um1dm2BaLntGLGYFmvKaOi8OU9EfZgdm8daPuUD16RVKsmHdSCWiZRFwluP5Lw5NRP0jnE5/KeNT
qnegFGpKdFMRu3Au17evtaMelATxdqBnkMG1zRSuWzEjdj1rwgs0+fUejl0CfuLnCuzsf2BpOS9s
bNAZcg0pkSSUbNcMmAqX66FURiAOg6ExzHCbyvJKFeNduNPrrERhWAqigTCX9TXFyZPtmjZLCGtd
ADpamrvSsM/6Z/Hluj6apC6qbey2+fNVop57R8YN5Oim8FIEEsQ1CPI6nra6evoSgYsbVop/voba
Y6EBygap6mgiSH2wzsAlTkM8V0X+PJX/eaPe1bIYnJvqDJ130L33hRlURCtkHKBgGixg7nt6XQpd
VHI6M6FehiqdA/8q0YQgke4LmFld3rOCIXfSgBQHiIP214yCRa+iZu0DAatVpTxTAG9UNcPVj6Kn
xJC6hV8XPPRN+4AnaBf13SMyYJ92n4O2jO5Rf2IB+N+i3UQh+4KlJAj67qu/dxXO4d7b0aUabPbi
QbsnzaVwSWdxHFHPMOVPBTMgg62lKOXBYHspK0w1UzQ73kkhQH43yl5mfcDskwRn18qxMsSRqqWz
IVeGtMRjJluwU0KMimBeMNxRG8UekwYLpjoMvk8Xr0Lp+T+zKAw1gCAwi0w4bidZC3UmDQu+psG9
+b3YwBXU6Mym2qItut7+vi/2xRge63EqueIXcDD0GdjAx3dlpA9ys6uin09iNwac/1v1hjjdPGbx
XEvIO9hwhvfqnc5/ZmB8pXNcndqFttsSdrpRg8+AYk4Y4prfivxbnhuLosJlnyXEWtr3zyZCOP7V
yRXb44Fozid5gCFTnlRTQStN1Vi8EAgnPpKfpBHpWpxTbg2LaVUEDZEXJwHIIQEABFj3vS+yPDXN
dPI5Qqiq2EhiwHrk1cpPmtfBgtqVBSu08wy1xyNaHgBEH5zMX9d4zY0Ji1oTq4TXVWVJj6pdlrrN
SU1AAHrX4snc/y14ZxPLqmPLsiQsHXjrV4l+YpTpVqsSee9p46NYdSELYx/0niEAfK5WWuBemqk+
45CJYe7Ko91+9EzI5kMhKLzjZPvfBjxwJy8zqqqBiVY4ZdUWZVgQRVHKIJkbn/wCBd5Ze1+cCDhh
JixperZCwn3BZW32VQLd8hOPjX8+bUIcDiNNR6fug6rovYzhpYjuiRLLW2RVBhsoUu3DWpOuy1g2
E9C2+wesKzClrhYowlyZhqH6T9/32MhQhfJxqgaTzjxYA53LGfPdO2RLVLviD/LNWqCii+UL2Bkl
E84aludCWMkJv9XEHcbD/XUf2ovwvAAbHHdbzMa3rnp2B6wos4eN0gohH23OZeGYJopeU2mTZQkN
dPqqClg7D29WRJsTwnHLZ9c8faKj5YcS2YZtl5x3iRXDA96TBDaymNnDPjW8uitIJWTGM78VKX8z
mZX5CLX29xw7EOqxDpWbJ5/bxUsvkXgMSxN+vbyld/DTArlbqpObn50LB0byWrlGvwcYLasTY5Xt
x4nU0b6hzGI2Gs6skH/Szw7OTXBng2yLvwu8adPsiVo5qWDTcfICDgCZd0R+c9Xc2yasPC+iHsvh
EtG5d9uLtzw89dHOxdxabOZkTzh/HCoX53eGznI6KugBa48OnsC4YE3DUsU+iafjlzI2YBDBlUrI
vQWRudwVF8dy0x3otobQGPsI4aCBqLe/ZLwPK/0lUqjqAwa+cEZUQlSHPpL+Y8dldAh6FHUKk1Y2
yKI3AkWcC58VXwFL37cnyad8q7kLMNOG2Vi7YL55ipI3ogVAMFL/aj3shL10sD8ryQUFaGkiPbUo
I2l0ettqiC5Acd8rgAN7yvGgvpvBoGFsOxJvQIeDKlItOElFRmY7lnUTZFq2e70yJM0J/J9xifkL
7DWO8ZOT/b4V9RoreuBLjb6Ad7fSV+xEMQu1hvnG4sUwfz7yC2JZvzZFEvi3iJDsZkxgRSgwrwFl
2QBfZneaJakq1g32p2H9OFHkYfc5FHA4mU8hizBbD6f5GYiVzDUpsVBquUU4/rWg34vMgNjUXdhy
3mdetSTfuFtydc3sJenQkTNW+WYYf1yubwtO2gIZMaQBNfttOss4qkI8lq91djHlH9i+VZ2PiMMj
+fBJkKuVOppSLGd88OK8PKaZ5tv0Soqu7JZyqM19IYRSRjJxhu4+0auFVxmT1ZTueQ93/WDxzumV
3VQnFhqdpllQ4q6AWf/M/hpT2+DN3d0zJoJT4t+pGnDu5idi47Wp0RieBPbLoEF6GYo0KxR5U+cN
JvduSM6FREGgUcEZ34hYj2Cx3LTwjn9ob9nIIiiHxitfKRRkJTUDsjTE/zcg2snvchdjuOJNxCbF
QZTPOHjrX/DL42XHI6BGbVINpfuhIlhExiLR1GSIlyi8QNMkRA7/cxrxkFPg+Pfs0Ex/vWP9RMQs
bxYdYUf1+VoUx4zQ9IowwkBiNi50BZcYjbHkY0+h0GYTesb9EHlJUKjuoQhy2NgXMyF3DsOy9ml0
CUu19a1uS1cW7bgPUh6CcFBhHzWrWgzihlFZmIGEjCQfmVF4zr+J177AGvzvWioAGkiT39q1a3B/
sX7vyOauDU9HkK7KDjg0Wc0raKaCFZ6Jw9GgVxMamZE/QUGAnq7K1C9zdZxmhdpVvJ35pcvkx5cL
sX01eEeTszp/+9TMxF96uScIdL7ua9kLBYv5L20WVzhBeDNXwkKv1S4BMVCUxLIbX+TbXinMGOOs
F0TMKzLJ0HSeeWEw9ol9mMYfBc9I/IC3+ekPUZiddtJi+DJvlIVxfZ+RuFiKct3O6z+AAqArDp7q
K6B5Fl3T8//qbLg9P2Lv7BQ2ItQZK/hlPUEDW7Hh95F/i4OAc2R9u4CYuctb5JpnhfE+g3HlR5Cm
WLAuXjfFpSDH2/Pp3Z9fp6bCCSJ/yJw4KxcYCdmGVnx9ljfkfh5ahVUCW+hIFHqIIOMGrv63RfkM
OuJkLO2MtlZ5GbVA/aIIGix3DhPSbp6LqqKV/02tcHN7FasI5J/GvB7mbWomdgxMDeJ8/5HhzZln
mepYziwzWSCorQocsNzVvevO4hMIVk1+a0XuMROAeE1Gf9vLEW4mUHl1USWnssjsAT6n0VCllDqg
/jxfPsebiQH3XmZm9OnY+U04eOzalu5AhlRrBpQxk8sNdrJVYAWr2lfAvoNd0h/40jmZLfcQeaLf
Xh+B/YD0LanpD0EqY5HSSaW61EAM+dVdKh26HhGM2bEQK0wmnGlbIzfeGzyNJ1BKJKUNMNGC8FiI
AH+1Z9K/IDGYu4vGH9Bmct6p3zdhUcB6rmX3tTC7IFAMMZSgYuISmIzy9NBRamB69hxhf4nxEt7/
ei40hxWnPiXtjwlonZKLJDZjV29RRtlnEbCHwiiecLBu5/k4bGZacoPP4wv6+sZMtmXraL/i4imG
GAnE6+8aCprON+xjSko9fHviOMSTGK50m9HAem7YSq4D3VailWnZY8nsnJ5fuueVQe4J0D6pMhUU
BS2cmlLl45KWP/xQUiiHH36u90b6tipd6sM8bnv6q54uDbabtHlGLn35LKcv0TblTxuwOol3p2rD
HzUXNIZZocmkLlJt0YUkotE35ZKVg41WOeH/HcBMQeqOMlZakke3OuybRViU2vkW26ivXry4QsuY
PSQIor6BLIAntYlY0aMZ1wXczw3G8UCEShiSgfBUDihIQ2mVg4BTANDiYb+F1RDuGAmMlLrmZRHe
mWUuT69vZ7nfLLJ0U28cx9Om/k4jKqIX6FVN4q2fhnNpTf57cgdE+xumuSey/recnTKZcHzzkREV
x+kL74TjEd1kcuONSVG4xMkat21tY7fbmklbESy2j+KUYzb3OAvxQ6AR7+G3nDWtITSFM18FqUv/
S+nSRD8wpuHQm42W4AkOuJh9OQkUoeKTfTfScmp39eG4NixkM870Lkr0CF3zRaLWNgDPjRAmP4E+
DOH9jKK1v9Ch04mna6iwvyIhzr8hqFoDmufShsRMyVKh032Epyg6XZxZrYN8C6FbKdbEWIDzlAQe
kPrAdUkwJ/p6MzFsGWZSRZ47hLOIvjwDzXgOMdKjJ0avH5L47worn11NBvyGcXf7nZ33Pc+c2JaO
VcM9xG4KTTf7+9rKUyQIABeaLT/nbYiO5N3Im6Q3kjf7L7ex0GZ/XRMsDGr8GMpc29oNf49x2QVt
laIT8lzrgAaDCdimkErD1UriEVhXxffFVH9rq5zTvkS7a+VSLKz3NerKtGsayoAHeGZHN/UNGju3
wAb4G6tsiI0t9dtn7qeedMOqoQdYVNa82T/b+WXh8PD8Vo5Po34fxEPurPgMSGNxvlsdOJAqkoTG
04yXxOgezVRS3m4lU8au+Wcg8uCl7f7UOKviRsQg/6WIcwzJWuNuv2kttqR3QTCMHDSuGc4pNKlh
6V0RStDlm6E3xM9nV0RNzPF9Qexxx0oTEcCTXsAGeoeyxIQtfhrH7GhOJtRCPCjhJ3XOejIm3a+y
H91wh1pGe+aQpwHP2cNpgD4rlPq8PWIVPovdLksvrkGg3cTqyG4QjMufhLdqHQ4izkAtVtYmmw8A
JndTW7UPetdVkXPX9kdLXj9hMiwPhadTVeW1iHmji2kb0Mn+31qQXkZ3tOFHv7HVuIRjOkwnroNs
JdqzWL2IBg7eP+ci1qe48WGP9HagNOQQ2vWI852Hu2nUplM1fAA7vXupj1+jX4nSqM1fKnSkN08X
k1CuclCC58XyCb0ZnHxBaHOWHQKxwuZThPHbE1VqWb5RgN4JvF5TpbZohSni9zqzoWZUI7bjjbzg
8s0uTuGL3jLgttmQUeQT1cvTBIup92SNq0YlQIDGF9lNrSclJ5ZTpmFhw3PAXXetr5C0z+8WZ4Wt
6eM/QMb+WvYtWQlHfAuQDpcUSjUva1JPfw5ZSuWrdazeV0mOBQCmaGXMleNGtrPdq7RoyBIA5NcA
Q/FDtgimNkkFjHyIelQ4z+t/Xc8atEzCLnuUs8bJHRQgWlhGD1M1VLV6BGZwDv0Y9CcP/yj3xk4l
t7GaTRdKc2VXouMjmHqZYWMDnwDyNfzYZ//OULp8YJuueqNfIiamhnkZ3gZ0GTLPWNnyIRv/EwXM
bj36B9Frty6rgIJ/AUvzpNKnvODqJT+DK3iLnlx+QzLiVDsT7Objm/qqyltmWaNt4+tvHw72HV2e
yQSyF1ZISb2HdkFtf7LJcdHy3nHz5m8MKlUv75j+PLbi3iyJrPGMZO6+/YIkLCNRVHNWOZCv/MUt
RV061NzdVoB+4XmPM381hPhHxq4pOWv/GICDb+kG4+9MZmb8jaKF+Zpq/zyypUcZb1lpwS6dXD8A
kFWMCmUJK26OBe/eMM34praqeBKTEr8fUukU1cuT0Vt6tyQZ1lyNwtiH0HjGGo9IydEcn3GLJd4g
jbq2I2zmAqTKhDA2dK/+ZRESmN0jn8fNbPSVavGNil71DYjno6yz
`protect end_protected
