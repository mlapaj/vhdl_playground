library IEEE;
use ieee.std_logic_1164.all;

entity top_module is
port (
   CLK: in std_logic
     );
end top_module;

architecture basic of top_module is

begin

end basic;